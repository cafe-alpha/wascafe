-- wasca.vhd

-- Generated using ACDS version 15.1 193

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity wasca is
	port (
		abus_slave_0_abus_address                      : in    std_logic_vector(9 downto 0)  := (others => '0'); --                 abus_slave_0_abus.address
		abus_slave_0_abus_chipselect                   : in    std_logic_vector(2 downto 0)  := (others => '0'); --                                  .chipselect
		abus_slave_0_abus_read                         : in    std_logic                     := '0';             --                                  .read
		abus_slave_0_abus_write                        : in    std_logic_vector(1 downto 0)  := (others => '0'); --                                  .write
		abus_slave_0_abus_waitrequest                  : out   std_logic;                                        --                                  .waitrequest
		abus_slave_0_abus_interrupt                    : out   std_logic;                                        --                                  .interrupt
		abus_slave_0_abus_addressdata                  : inout std_logic_vector(15 downto 0) := (others => '0'); --                                  .addressdata
		abus_slave_0_abus_direction                    : out   std_logic;                                        --                                  .direction
		abus_slave_0_abus_muxing                       : out   std_logic_vector(1 downto 0);                     --                                  .muxing
		abus_slave_0_abus_disableout                   : out   std_logic;                                        --                                  .disableout
		abus_slave_0_conduit_saturn_reset_saturn_reset : in    std_logic                     := '0';             -- abus_slave_0_conduit_saturn_reset.saturn_reset
		altpll_0_areset_conduit_export                 : in    std_logic                     := '0';             --           altpll_0_areset_conduit.export
		altpll_0_locked_conduit_export                 : out   std_logic;                                        --           altpll_0_locked_conduit.export
		altpll_0_phasedone_conduit_export              : out   std_logic;                                        --        altpll_0_phasedone_conduit.export
		clk_clk                                        : in    std_logic                     := '0';             --                               clk.clk
		clock_116_mhz_clk                              : out   std_logic;                                        --                     clock_116_mhz.clk
		external_sdram_controller_wire_addr            : out   std_logic_vector(12 downto 0);                    --    external_sdram_controller_wire.addr
		external_sdram_controller_wire_ba              : out   std_logic_vector(1 downto 0);                     --                                  .ba
		external_sdram_controller_wire_cas_n           : out   std_logic;                                        --                                  .cas_n
		external_sdram_controller_wire_cke             : out   std_logic;                                        --                                  .cke
		external_sdram_controller_wire_cs_n            : out   std_logic;                                        --                                  .cs_n
		external_sdram_controller_wire_dq              : inout std_logic_vector(15 downto 0) := (others => '0'); --                                  .dq
		external_sdram_controller_wire_dqm             : out   std_logic_vector(1 downto 0);                     --                                  .dqm
		external_sdram_controller_wire_ras_n           : out   std_logic;                                        --                                  .ras_n
		external_sdram_controller_wire_we_n            : out   std_logic;                                        --                                  .we_n
		leds_conn_export                               : out   std_logic_vector(3 downto 0);                     --                         leds_conn.export
		sdram_clkout_clk                               : out   std_logic;                                        --                      sdram_clkout.clk
		switches_conn_export                           : in    std_logic_vector(2 downto 0)  := (others => '0'); --                     switches_conn.export
		uart_0_external_connection_rxd                 : in    std_logic                     := '0';             --        uart_0_external_connection.rxd
		uart_0_external_connection_txd                 : out   std_logic                                         --                                  .txd
	);
end entity wasca;

architecture rtl of wasca is
	component abus_demux is
		port (
			clock                     : in    std_logic                     := 'X';             -- clk
			abus_address              : in    std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			abus_chipselect           : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- chipselect
			abus_read                 : in    std_logic                     := 'X';             -- read
			abus_write                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- write
			abus_waitrequest          : out   std_logic;                                        -- waitrequest
			abus_interrupt            : out   std_logic;                                        -- interrupt
			abus_addressdata          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- addressdata
			abus_direction            : out   std_logic;                                        -- direction
			abus_muxing               : out   std_logic_vector(1 downto 0);                     -- muxing
			abus_disable_out          : out   std_logic;                                        -- disableout
			reset                     : in    std_logic                     := 'X';             -- reset
			avalon_nios_read          : in    std_logic                     := 'X';             -- read
			avalon_nios_write         : in    std_logic                     := 'X';             -- write
			avalon_nios_address       : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avalon_nios_writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avalon_nios_readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			avalon_nios_waitrequest   : out   std_logic;                                        -- waitrequest
			avalon_nios_readdatavalid : out   std_logic;                                        -- readdatavalid
			avalon_nios_burstcount    : in    std_logic                     := 'X';             -- burstcount
			demux_writeaddress        : out   std_logic_vector(27 downto 0);                    -- writeaddress
			demux_writedata           : out   std_logic_vector(15 downto 0);                    -- data
			demux_writepulse          : out   std_logic;                                        -- writepulse
			demux_write_byteenable    : out   std_logic_vector(1 downto 0);                     -- write_byteenable
			demux_readdata            : in    std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			demux_readpulse           : out   std_logic;                                        -- readpulse
			demux_readdatavalid       : in    std_logic                     := 'X';             -- readdatavalid
			demux_readaddress         : out   std_logic_vector(27 downto 0);                    -- readaddress
			saturn_reset              : in    std_logic                     := 'X'              -- saturn_reset
		);
	end component abus_demux;

	component abus_slave is
		port (
			clock                     : in  std_logic                     := 'X';             -- clk
			avalon_read               : out std_logic;                                        -- read
			avalon_write              : out std_logic;                                        -- write
			avalon_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			avalon_address            : out std_logic_vector(27 downto 0);                    -- address
			avalon_readdata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			avalon_writedata          : out std_logic_vector(15 downto 0);                    -- writedata
			avalon_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			avalon_burstcount         : out std_logic;                                        -- burstcount
			reset                     : in  std_logic                     := 'X';             -- reset
			avalon_nios_read          : in  std_logic                     := 'X';             -- read
			avalon_nios_write         : in  std_logic                     := 'X';             -- write
			avalon_nios_address       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avalon_nios_writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avalon_nios_readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			avalon_nios_waitrequest   : out std_logic;                                        -- waitrequest
			avalon_nios_readdatavalid : out std_logic;                                        -- readdatavalid
			avalon_nios_burstcount    : in  std_logic                     := 'X';             -- burstcount
			demux_writeaddress        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- writeaddress
			demux_writedata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			demux_writepulse          : in  std_logic                     := 'X';             -- writepulse
			demux_write_byteenable    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- write_byteenable
			demux_readdata            : out std_logic_vector(15 downto 0);                    -- readdata
			demux_readpulse           : in  std_logic                     := 'X';             -- readpulse
			demux_readdatavalid       : out std_logic;                                        -- readdatavalid
			demux_readaddress         : in  std_logic_vector(27 downto 0) := (others => 'X')  -- readaddress
		);
	end component abus_slave;

	component wasca_altpll_0 is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			c1        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component wasca_altpll_0;

	component wasca_external_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component wasca_external_sdram_controller;

	component wasca_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component wasca_leds;

	component wasca_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component wasca_nios2_gen2_0;

	component altera_onchip_flash is
		generic (
			INIT_FILENAME                       : string  := "";
			INIT_FILENAME_SIM                   : string  := "";
			DEVICE_FAMILY                       : string  := "Unknown";
			PART_NAME                           : string  := "Unknown";
			DEVICE_ID                           : string  := "Unknown";
			SECTOR1_START_ADDR                  : integer := 0;
			SECTOR1_END_ADDR                    : integer := 0;
			SECTOR2_START_ADDR                  : integer := 0;
			SECTOR2_END_ADDR                    : integer := 0;
			SECTOR3_START_ADDR                  : integer := 0;
			SECTOR3_END_ADDR                    : integer := 0;
			SECTOR4_START_ADDR                  : integer := 0;
			SECTOR4_END_ADDR                    : integer := 0;
			SECTOR5_START_ADDR                  : integer := 0;
			SECTOR5_END_ADDR                    : integer := 0;
			MIN_VALID_ADDR                      : integer := 0;
			MAX_VALID_ADDR                      : integer := 0;
			MIN_UFM_VALID_ADDR                  : integer := 0;
			MAX_UFM_VALID_ADDR                  : integer := 0;
			SECTOR1_MAP                         : integer := 0;
			SECTOR2_MAP                         : integer := 0;
			SECTOR3_MAP                         : integer := 0;
			SECTOR4_MAP                         : integer := 0;
			SECTOR5_MAP                         : integer := 0;
			ADDR_RANGE1_END_ADDR                : integer := 0;
			ADDR_RANGE1_OFFSET                  : integer := 0;
			ADDR_RANGE2_OFFSET                  : integer := 0;
			AVMM_DATA_ADDR_WIDTH                : integer := 19;
			AVMM_DATA_DATA_WIDTH                : integer := 32;
			AVMM_DATA_BURSTCOUNT_WIDTH          : integer := 4;
			SECTOR_READ_PROTECTION_MODE         : integer := 31;
			FLASH_SEQ_READ_DATA_COUNT           : integer := 2;
			FLASH_ADDR_ALIGNMENT_BITS           : integer := 1;
			FLASH_READ_CYCLE_MAX_INDEX          : integer := 4;
			FLASH_RESET_CYCLE_MAX_INDEX         : integer := 29;
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  : integer := 112;
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX : integer := 40603248;
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX : integer := 35382;
			PARALLEL_MODE                       : boolean := true;
			READ_AND_WRITE_MODE                 : boolean := true;
			WRAPPING_BURST_MODE                 : boolean := false;
			IS_DUAL_BOOT                        : string  := "False";
			IS_ERAM_SKIP                        : string  := "False";
			IS_COMPRESSED_IMAGE                 : string  := "False"
		);
		port (
			clock                   : in  std_logic                     := 'X';             -- clk
			reset_n                 : in  std_logic                     := 'X';             -- reset_n
			avmm_data_addr          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			avmm_data_read          : in  std_logic                     := 'X';             -- read
			avmm_data_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_data_write         : in  std_logic                     := 'X';             -- write
			avmm_data_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_data_waitrequest   : out std_logic;                                        -- waitrequest
			avmm_data_readdatavalid : out std_logic;                                        -- readdatavalid
			avmm_data_burstcount    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			avmm_csr_addr           : in  std_logic                     := 'X';             -- address
			avmm_csr_read           : in  std_logic                     := 'X';             -- read
			avmm_csr_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_csr_write          : in  std_logic                     := 'X';             -- write
			avmm_csr_readdata       : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_onchip_flash;

	component wasca_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component wasca_onchip_memory2_0;

	component wasca_onchip_memory2_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component wasca_onchip_memory2_1;

	component wasca_performance_counter_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component wasca_performance_counter_0;

	component wasca_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- export
		);
	end component wasca_switches;

	component wasca_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			dataavailable : out std_logic;                                        -- dataavailable
			readyfordata  : out std_logic;                                        -- readyfordata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component wasca_uart_0;

	component wasca_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                              : in  std_logic                     := 'X';             -- clk
			abus_slave_0_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			abus_slave_0_avalon_master_address                         : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			abus_slave_0_avalon_master_waitrequest                     : out std_logic;                                        -- waitrequest
			abus_slave_0_avalon_master_burstcount                      : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			abus_slave_0_avalon_master_read                            : in  std_logic                     := 'X';             -- read
			abus_slave_0_avalon_master_readdata                        : out std_logic_vector(15 downto 0);                    -- readdata
			abus_slave_0_avalon_master_readdatavalid                   : out std_logic;                                        -- readdatavalid
			abus_slave_0_avalon_master_write                           : in  std_logic                     := 'X';             -- write
			abus_slave_0_avalon_master_writedata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_address                           : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                       : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                              : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                             : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                    : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                       : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			abus_demux_0_avalon_nios_address                           : out std_logic_vector(7 downto 0);                     -- address
			abus_demux_0_avalon_nios_write                             : out std_logic;                                        -- write
			abus_demux_0_avalon_nios_read                              : out std_logic;                                        -- read
			abus_demux_0_avalon_nios_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			abus_demux_0_avalon_nios_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			abus_demux_0_avalon_nios_burstcount                        : out std_logic_vector(0 downto 0);                     -- burstcount
			abus_demux_0_avalon_nios_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			abus_demux_0_avalon_nios_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			abus_slave_0_avalon_nios_address                           : out std_logic_vector(7 downto 0);                     -- address
			abus_slave_0_avalon_nios_write                             : out std_logic;                                        -- write
			abus_slave_0_avalon_nios_read                              : out std_logic;                                        -- read
			abus_slave_0_avalon_nios_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			abus_slave_0_avalon_nios_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			abus_slave_0_avalon_nios_burstcount                        : out std_logic_vector(0 downto 0);                     -- burstcount
			abus_slave_0_avalon_nios_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			abus_slave_0_avalon_nios_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			altpll_0_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                   : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                    : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			external_sdram_controller_s1_address                       : out std_logic_vector(23 downto 0);                    -- address
			external_sdram_controller_s1_write                         : out std_logic;                                        -- write
			external_sdram_controller_s1_read                          : out std_logic;                                        -- read
			external_sdram_controller_s1_readdata                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			external_sdram_controller_s1_writedata                     : out std_logic_vector(15 downto 0);                    -- writedata
			external_sdram_controller_s1_byteenable                    : out std_logic_vector(1 downto 0);                     -- byteenable
			external_sdram_controller_s1_readdatavalid                 : in  std_logic                     := 'X';             -- readdatavalid
			external_sdram_controller_s1_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			external_sdram_controller_s1_chipselect                    : out std_logic;                                        -- chipselect
			leds_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                              : out std_logic;                                        -- write
			leds_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                                         : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                       : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                         : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                          : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                   : out std_logic;                                        -- debugaccess
			onchip_flash_0_csr_address                                 : out std_logic_vector(0 downto 0);                     -- address
			onchip_flash_0_csr_write                                   : out std_logic;                                        -- write
			onchip_flash_0_csr_read                                    : out std_logic;                                        -- read
			onchip_flash_0_csr_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_0_csr_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_0_data_address                                : out std_logic_vector(15 downto 0);                    -- address
			onchip_flash_0_data_write                                  : out std_logic;                                        -- write
			onchip_flash_0_data_read                                   : out std_logic;                                        -- read
			onchip_flash_0_data_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_0_data_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_0_data_burstcount                             : out std_logic_vector(3 downto 0);                     -- burstcount
			onchip_flash_0_data_readdatavalid                          : in  std_logic                     := 'X';             -- readdatavalid
			onchip_flash_0_data_waitrequest                            : in  std_logic                     := 'X';             -- waitrequest
			onchip_memory2_0_s1_address                                : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_0_s1_write                                  : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                  : out std_logic;                                        -- clken
			onchip_memory2_1_s1_address                                : out std_logic_vector(9 downto 0);                     -- address
			onchip_memory2_1_s1_write                                  : out std_logic;                                        -- write
			onchip_memory2_1_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_1_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_1_s1_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_1_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory2_1_s1_clken                                  : out std_logic;                                        -- clken
			performance_counter_0_control_slave_address                : out std_logic_vector(2 downto 0);                     -- address
			performance_counter_0_control_slave_write                  : out std_logic;                                        -- write
			performance_counter_0_control_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			performance_counter_0_control_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			performance_counter_0_control_slave_begintransfer          : out std_logic;                                        -- begintransfer
			switches_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_address                                          : out std_logic_vector(2 downto 0);                     -- address
			uart_0_s1_write                                            : out std_logic;                                        -- write
			uart_0_s1_read                                             : out std_logic;                                        -- read
			uart_0_s1_readdata                                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_writedata                                        : out std_logic_vector(15 downto 0);                    -- writedata
			uart_0_s1_begintransfer                                    : out std_logic;                                        -- begintransfer
			uart_0_s1_chipselect                                       : out std_logic                                         -- chipselect
		);
	end component wasca_mm_interconnect_0;

	component wasca_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component wasca_irq_mapper;

	component wasca_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component wasca_rst_controller;

	component wasca_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component wasca_rst_controller_001;

	signal altpll_0_c0_clk                                                     : std_logic;                     -- altpll_0:c0 -> [clock_116_mhz_clk, abus_demux_0:clock, abus_slave_0:clock, external_sdram_controller:clk, irq_mapper:clk, leds:clk, mm_interconnect_0:altpll_0_c0_clk, nios2_gen2_0:clk, onchip_flash_0:clock, onchip_memory2_0:clk, onchip_memory2_1:clk, performance_counter_0:clk, rst_controller:clk, rst_controller_002:clk, switches:clk, uart_0:clk]
	signal abus_slave_0_demux_readdata                                         : std_logic_vector(15 downto 0); -- abus_slave_0:demux_readdata -> abus_demux_0:demux_readdata
	signal abus_demux_0_demux_readpulse                                        : std_logic;                     -- abus_demux_0:demux_readpulse -> abus_slave_0:demux_readpulse
	signal abus_demux_0_demux_readaddress                                      : std_logic_vector(27 downto 0); -- abus_demux_0:demux_readaddress -> abus_slave_0:demux_readaddress
	signal abus_demux_0_demux_data                                             : std_logic_vector(15 downto 0); -- abus_demux_0:demux_writedata -> abus_slave_0:demux_writedata
	signal abus_slave_0_demux_readdatavalid                                    : std_logic;                     -- abus_slave_0:demux_readdatavalid -> abus_demux_0:demux_readdatavalid
	signal abus_demux_0_demux_write_byteenable                                 : std_logic_vector(1 downto 0);  -- abus_demux_0:demux_write_byteenable -> abus_slave_0:demux_write_byteenable
	signal abus_demux_0_demux_writeaddress                                     : std_logic_vector(27 downto 0); -- abus_demux_0:demux_writeaddress -> abus_slave_0:demux_writeaddress
	signal abus_demux_0_demux_writepulse                                       : std_logic;                     -- abus_demux_0:demux_writepulse -> abus_slave_0:demux_writepulse
	signal nios2_gen2_0_debug_reset_request_reset                              : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal abus_slave_0_avalon_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:abus_slave_0_avalon_master_waitrequest -> abus_slave_0:avalon_waitrequest
	signal abus_slave_0_avalon_master_readdata                                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:abus_slave_0_avalon_master_readdata -> abus_slave_0:avalon_readdata
	signal abus_slave_0_avalon_master_read                                     : std_logic;                     -- abus_slave_0:avalon_read -> mm_interconnect_0:abus_slave_0_avalon_master_read
	signal abus_slave_0_avalon_master_address                                  : std_logic_vector(27 downto 0); -- abus_slave_0:avalon_address -> mm_interconnect_0:abus_slave_0_avalon_master_address
	signal abus_slave_0_avalon_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:abus_slave_0_avalon_master_readdatavalid -> abus_slave_0:avalon_readdatavalid
	signal abus_slave_0_avalon_master_write                                    : std_logic;                     -- abus_slave_0:avalon_write -> mm_interconnect_0:abus_slave_0_avalon_master_write
	signal abus_slave_0_avalon_master_writedata                                : std_logic_vector(15 downto 0); -- abus_slave_0:avalon_writedata -> mm_interconnect_0:abus_slave_0_avalon_master_writedata
	signal abus_slave_0_avalon_master_burstcount                               : std_logic;                     -- abus_slave_0:avalon_burstcount -> mm_interconnect_0:abus_slave_0_avalon_master_burstcount
	signal nios2_gen2_0_data_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                    : std_logic_vector(26 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                 : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                       : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                      : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                  : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                             : std_logic_vector(26 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_external_sdram_controller_s1_chipselect           : std_logic;                     -- mm_interconnect_0:external_sdram_controller_s1_chipselect -> external_sdram_controller:az_cs
	signal mm_interconnect_0_external_sdram_controller_s1_readdata             : std_logic_vector(15 downto 0); -- external_sdram_controller:za_data -> mm_interconnect_0:external_sdram_controller_s1_readdata
	signal mm_interconnect_0_external_sdram_controller_s1_waitrequest          : std_logic;                     -- external_sdram_controller:za_waitrequest -> mm_interconnect_0:external_sdram_controller_s1_waitrequest
	signal mm_interconnect_0_external_sdram_controller_s1_address              : std_logic_vector(23 downto 0); -- mm_interconnect_0:external_sdram_controller_s1_address -> external_sdram_controller:az_addr
	signal mm_interconnect_0_external_sdram_controller_s1_read                 : std_logic;                     -- mm_interconnect_0:external_sdram_controller_s1_read -> mm_interconnect_0_external_sdram_controller_s1_read:in
	signal mm_interconnect_0_external_sdram_controller_s1_byteenable           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:external_sdram_controller_s1_byteenable -> mm_interconnect_0_external_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_external_sdram_controller_s1_readdatavalid        : std_logic;                     -- external_sdram_controller:za_valid -> mm_interconnect_0:external_sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_external_sdram_controller_s1_write                : std_logic;                     -- mm_interconnect_0:external_sdram_controller_s1_write -> mm_interconnect_0_external_sdram_controller_s1_write:in
	signal mm_interconnect_0_external_sdram_controller_s1_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_0:external_sdram_controller_s1_writedata -> external_sdram_controller:az_data
	signal mm_interconnect_0_onchip_memory2_1_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	signal mm_interconnect_0_onchip_memory2_1_s1_readdata                      : std_logic_vector(31 downto 0); -- onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	signal mm_interconnect_0_onchip_memory2_1_s1_address                       : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	signal mm_interconnect_0_onchip_memory2_1_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	signal mm_interconnect_0_onchip_memory2_1_s1_write                         : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	signal mm_interconnect_0_onchip_memory2_1_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	signal mm_interconnect_0_onchip_memory2_1_s1_clken                         : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	signal mm_interconnect_0_abus_slave_0_avalon_nios_readdata                 : std_logic_vector(15 downto 0); -- abus_slave_0:avalon_nios_readdata -> mm_interconnect_0:abus_slave_0_avalon_nios_readdata
	signal mm_interconnect_0_abus_slave_0_avalon_nios_waitrequest              : std_logic;                     -- abus_slave_0:avalon_nios_waitrequest -> mm_interconnect_0:abus_slave_0_avalon_nios_waitrequest
	signal mm_interconnect_0_abus_slave_0_avalon_nios_address                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:abus_slave_0_avalon_nios_address -> abus_slave_0:avalon_nios_address
	signal mm_interconnect_0_abus_slave_0_avalon_nios_read                     : std_logic;                     -- mm_interconnect_0:abus_slave_0_avalon_nios_read -> abus_slave_0:avalon_nios_read
	signal mm_interconnect_0_abus_slave_0_avalon_nios_readdatavalid            : std_logic;                     -- abus_slave_0:avalon_nios_readdatavalid -> mm_interconnect_0:abus_slave_0_avalon_nios_readdatavalid
	signal mm_interconnect_0_abus_slave_0_avalon_nios_write                    : std_logic;                     -- mm_interconnect_0:abus_slave_0_avalon_nios_write -> abus_slave_0:avalon_nios_write
	signal mm_interconnect_0_abus_slave_0_avalon_nios_writedata                : std_logic_vector(15 downto 0); -- mm_interconnect_0:abus_slave_0_avalon_nios_writedata -> abus_slave_0:avalon_nios_writedata
	signal mm_interconnect_0_abus_slave_0_avalon_nios_burstcount               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:abus_slave_0_avalon_nios_burstcount -> abus_slave_0:avalon_nios_burstcount
	signal mm_interconnect_0_abus_demux_0_avalon_nios_readdata                 : std_logic_vector(15 downto 0); -- abus_demux_0:avalon_nios_readdata -> mm_interconnect_0:abus_demux_0_avalon_nios_readdata
	signal mm_interconnect_0_abus_demux_0_avalon_nios_waitrequest              : std_logic;                     -- abus_demux_0:avalon_nios_waitrequest -> mm_interconnect_0:abus_demux_0_avalon_nios_waitrequest
	signal mm_interconnect_0_abus_demux_0_avalon_nios_address                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:abus_demux_0_avalon_nios_address -> abus_demux_0:avalon_nios_address
	signal mm_interconnect_0_abus_demux_0_avalon_nios_read                     : std_logic;                     -- mm_interconnect_0:abus_demux_0_avalon_nios_read -> abus_demux_0:avalon_nios_read
	signal mm_interconnect_0_abus_demux_0_avalon_nios_readdatavalid            : std_logic;                     -- abus_demux_0:avalon_nios_readdatavalid -> mm_interconnect_0:abus_demux_0_avalon_nios_readdatavalid
	signal mm_interconnect_0_abus_demux_0_avalon_nios_write                    : std_logic;                     -- mm_interconnect_0:abus_demux_0_avalon_nios_write -> abus_demux_0:avalon_nios_write
	signal mm_interconnect_0_abus_demux_0_avalon_nios_writedata                : std_logic_vector(15 downto 0); -- mm_interconnect_0:abus_demux_0_avalon_nios_writedata -> abus_demux_0:avalon_nios_writedata
	signal mm_interconnect_0_abus_demux_0_avalon_nios_burstcount               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:abus_demux_0_avalon_nios_burstcount -> abus_demux_0:avalon_nios_burstcount
	signal mm_interconnect_0_onchip_flash_0_csr_readdata                       : std_logic_vector(31 downto 0); -- onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	signal mm_interconnect_0_onchip_flash_0_csr_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	signal mm_interconnect_0_onchip_flash_0_csr_read                           : std_logic;                     -- mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	signal mm_interconnect_0_onchip_flash_0_csr_write                          : std_logic;                     -- mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	signal mm_interconnect_0_onchip_flash_0_csr_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	signal mm_interconnect_0_onchip_flash_0_data_readdata                      : std_logic_vector(31 downto 0); -- onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	signal mm_interconnect_0_onchip_flash_0_data_waitrequest                   : std_logic;                     -- onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	signal mm_interconnect_0_onchip_flash_0_data_address                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	signal mm_interconnect_0_onchip_flash_0_data_read                          : std_logic;                     -- mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	signal mm_interconnect_0_onchip_flash_0_data_readdatavalid                 : std_logic;                     -- onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	signal mm_interconnect_0_onchip_flash_0_data_write                         : std_logic;                     -- mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	signal mm_interconnect_0_onchip_flash_0_data_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	signal mm_interconnect_0_onchip_flash_0_data_burstcount                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata             : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest          : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address              : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                 : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                      : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                       : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                         : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                         : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_performance_counter_0_control_slave_readdata      : std_logic_vector(31 downto 0); -- performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	signal mm_interconnect_0_performance_counter_0_control_slave_address       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	signal mm_interconnect_0_performance_counter_0_control_slave_begintransfer : std_logic;                     -- mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	signal mm_interconnect_0_performance_counter_0_control_slave_write         : std_logic;                     -- mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	signal mm_interconnect_0_performance_counter_0_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                       : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                           : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                          : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_switches_s1_readdata                              : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal mm_interconnect_0_leds_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                                  : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                                     : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_uart_0_s1_chipselect                              : std_logic;                     -- mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	signal mm_interconnect_0_uart_0_s1_readdata                                : std_logic_vector(15 downto 0); -- uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	signal mm_interconnect_0_uart_0_s1_address                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_0_s1_address -> uart_0:address
	signal mm_interconnect_0_uart_0_s1_read                                    : std_logic;                     -- mm_interconnect_0:uart_0_s1_read -> mm_interconnect_0_uart_0_s1_read:in
	signal mm_interconnect_0_uart_0_s1_begintransfer                           : std_logic;                     -- mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	signal mm_interconnect_0_uart_0_s1_write                                   : std_logic;                     -- mm_interconnect_0:uart_0_s1_write -> mm_interconnect_0_uart_0_s1_write:in
	signal mm_interconnect_0_uart_0_s1_writedata                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- uart_0:irq -> irq_mapper:receiver0_irq
	signal nios2_gen2_0_irq_irq                                                : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [abus_demux_0:reset, abus_slave_0:reset, irq_mapper:reset, mm_interconnect_0:abus_slave_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, onchip_memory2_1:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                  : std_logic;                     -- rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_1:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	signal mm_interconnect_0_external_sdram_controller_s1_read_ports_inv       : std_logic;                     -- mm_interconnect_0_external_sdram_controller_s1_read:inv -> external_sdram_controller:az_rd_n
	signal mm_interconnect_0_external_sdram_controller_s1_byteenable_ports_inv : std_logic_vector(1 downto 0);  -- mm_interconnect_0_external_sdram_controller_s1_byteenable:inv -> external_sdram_controller:az_be_n
	signal mm_interconnect_0_external_sdram_controller_s1_write_ports_inv      : std_logic;                     -- mm_interconnect_0_external_sdram_controller_s1_write:inv -> external_sdram_controller:az_wr_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal mm_interconnect_0_uart_0_s1_read_ports_inv                          : std_logic;                     -- mm_interconnect_0_uart_0_s1_read:inv -> uart_0:read_n
	signal mm_interconnect_0_uart_0_s1_write_ports_inv                         : std_logic;                     -- mm_interconnect_0_uart_0_s1_write:inv -> uart_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [external_sdram_controller:reset_n, leds:reset_n, nios2_gen2_0:reset_n, onchip_flash_0:reset_n, performance_counter_0:reset_n, switches:reset_n, uart_0:reset_n]

begin

	abus_demux_0 : component abus_demux
		port map (
			clock                     => altpll_0_c0_clk,                                          --                clock.clk
			abus_address              => abus_slave_0_abus_address,                                --                 abus.address
			abus_chipselect           => abus_slave_0_abus_chipselect,                             --                     .chipselect
			abus_read                 => abus_slave_0_abus_read,                                   --                     .read
			abus_write                => abus_slave_0_abus_write,                                  --                     .write
			abus_waitrequest          => abus_slave_0_abus_waitrequest,                            --                     .waitrequest
			abus_interrupt            => abus_slave_0_abus_interrupt,                              --                     .interrupt
			abus_addressdata          => abus_slave_0_abus_addressdata,                            --                     .addressdata
			abus_direction            => abus_slave_0_abus_direction,                              --                     .direction
			abus_muxing               => abus_slave_0_abus_muxing,                                 --                     .muxing
			abus_disable_out          => abus_slave_0_abus_disableout,                             --                     .disableout
			reset                     => rst_controller_reset_out_reset,                           --                reset.reset
			avalon_nios_read          => mm_interconnect_0_abus_demux_0_avalon_nios_read,          --          avalon_nios.read
			avalon_nios_write         => mm_interconnect_0_abus_demux_0_avalon_nios_write,         --                     .write
			avalon_nios_address       => mm_interconnect_0_abus_demux_0_avalon_nios_address,       --                     .address
			avalon_nios_writedata     => mm_interconnect_0_abus_demux_0_avalon_nios_writedata,     --                     .writedata
			avalon_nios_readdata      => mm_interconnect_0_abus_demux_0_avalon_nios_readdata,      --                     .readdata
			avalon_nios_waitrequest   => mm_interconnect_0_abus_demux_0_avalon_nios_waitrequest,   --                     .waitrequest
			avalon_nios_readdatavalid => mm_interconnect_0_abus_demux_0_avalon_nios_readdatavalid, --                     .readdatavalid
			avalon_nios_burstcount    => mm_interconnect_0_abus_demux_0_avalon_nios_burstcount(0), --                     .burstcount
			demux_writeaddress        => abus_demux_0_demux_writeaddress,                          --                demux.writeaddress
			demux_writedata           => abus_demux_0_demux_data,                                  --                     .data
			demux_writepulse          => abus_demux_0_demux_writepulse,                            --                     .writepulse
			demux_write_byteenable    => abus_demux_0_demux_write_byteenable,                      --                     .write_byteenable
			demux_readdata            => abus_slave_0_demux_readdata,                              --                     .readdata
			demux_readpulse           => abus_demux_0_demux_readpulse,                             --                     .readpulse
			demux_readdatavalid       => abus_slave_0_demux_readdatavalid,                         --                     .readdatavalid
			demux_readaddress         => abus_demux_0_demux_readaddress,                           --                     .readaddress
			saturn_reset              => abus_slave_0_conduit_saturn_reset_saturn_reset            -- conduit_saturn_reset.saturn_reset
		);

	abus_slave_0 : component abus_slave
		port map (
			clock                     => altpll_0_c0_clk,                                          --         clock.clk
			avalon_read               => abus_slave_0_avalon_master_read,                          -- avalon_master.read
			avalon_write              => abus_slave_0_avalon_master_write,                         --              .write
			avalon_waitrequest        => abus_slave_0_avalon_master_waitrequest,                   --              .waitrequest
			avalon_address            => abus_slave_0_avalon_master_address,                       --              .address
			avalon_readdata           => abus_slave_0_avalon_master_readdata,                      --              .readdata
			avalon_writedata          => abus_slave_0_avalon_master_writedata,                     --              .writedata
			avalon_readdatavalid      => abus_slave_0_avalon_master_readdatavalid,                 --              .readdatavalid
			avalon_burstcount         => abus_slave_0_avalon_master_burstcount,                    --              .burstcount
			reset                     => rst_controller_reset_out_reset,                           --         reset.reset
			avalon_nios_read          => mm_interconnect_0_abus_slave_0_avalon_nios_read,          --   avalon_nios.read
			avalon_nios_write         => mm_interconnect_0_abus_slave_0_avalon_nios_write,         --              .write
			avalon_nios_address       => mm_interconnect_0_abus_slave_0_avalon_nios_address,       --              .address
			avalon_nios_writedata     => mm_interconnect_0_abus_slave_0_avalon_nios_writedata,     --              .writedata
			avalon_nios_readdata      => mm_interconnect_0_abus_slave_0_avalon_nios_readdata,      --              .readdata
			avalon_nios_waitrequest   => mm_interconnect_0_abus_slave_0_avalon_nios_waitrequest,   --              .waitrequest
			avalon_nios_readdatavalid => mm_interconnect_0_abus_slave_0_avalon_nios_readdatavalid, --              .readdatavalid
			avalon_nios_burstcount    => mm_interconnect_0_abus_slave_0_avalon_nios_burstcount(0), --              .burstcount
			demux_writeaddress        => abus_demux_0_demux_writeaddress,                          --         demux.writeaddress
			demux_writedata           => abus_demux_0_demux_data,                                  --              .data
			demux_writepulse          => abus_demux_0_demux_writepulse,                            --              .writepulse
			demux_write_byteenable    => abus_demux_0_demux_write_byteenable,                      --              .write_byteenable
			demux_readdata            => abus_slave_0_demux_readdata,                              --              .readdata
			demux_readpulse           => abus_demux_0_demux_readpulse,                             --              .readpulse
			demux_readdatavalid       => abus_slave_0_demux_readdatavalid,                         --              .readdatavalid
			demux_readaddress         => abus_demux_0_demux_readaddress                            --              .readaddress
		);

	altpll_0 : component wasca_altpll_0
		port map (
			clk       => clk_clk,                                        --       inclk_interface.clk
			reset     => rst_controller_001_reset_out_reset,             -- inclk_interface_reset.reset
			read      => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write     => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address   => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata  => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0        => altpll_0_c0_clk,                                --                    c0.clk
			c1        => sdram_clkout_clk,                               --                    c1.clk
			areset    => altpll_0_areset_conduit_export,                 --        areset_conduit.export
			locked    => altpll_0_locked_conduit_export,                 --        locked_conduit.export
			phasedone => altpll_0_phasedone_conduit_export               --     phasedone_conduit.export
		);

	external_sdram_controller : component wasca_external_sdram_controller
		port map (
			clk            => altpll_0_c0_clk,                                                     --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                            -- reset.reset_n
			az_addr        => mm_interconnect_0_external_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_external_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_external_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_external_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_external_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_external_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_external_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_external_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_external_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => external_sdram_controller_wire_addr,                                 --  wire.export
			zs_ba          => external_sdram_controller_wire_ba,                                   --      .export
			zs_cas_n       => external_sdram_controller_wire_cas_n,                                --      .export
			zs_cke         => external_sdram_controller_wire_cke,                                  --      .export
			zs_cs_n        => external_sdram_controller_wire_cs_n,                                 --      .export
			zs_dq          => external_sdram_controller_wire_dq,                                   --      .export
			zs_dqm         => external_sdram_controller_wire_dqm,                                  --      .export
			zs_ras_n       => external_sdram_controller_wire_ras_n,                                --      .export
			zs_we_n        => external_sdram_controller_wire_we_n                                  --      .export
		);

	leds : component wasca_leds
		port map (
			clk        => altpll_0_c0_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_conn_export                           -- external_connection.export
		);

	nios2_gen2_0 : component wasca_nios2_gen2_0
		port map (
			clk                                 => altpll_0_c0_clk,                                            --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_flash_0 : component altera_onchip_flash
		generic map (
			INIT_FILENAME                       => "",
			INIT_FILENAME_SIM                   => "",
			DEVICE_FAMILY                       => "MAX 10",
			PART_NAME                           => "10M08SCE144C8G",
			DEVICE_ID                           => "08",
			SECTOR1_START_ADDR                  => 0,
			SECTOR1_END_ADDR                    => 4095,
			SECTOR2_START_ADDR                  => 4096,
			SECTOR2_END_ADDR                    => 8191,
			SECTOR3_START_ADDR                  => 8192,
			SECTOR3_END_ADDR                    => 23039,
			SECTOR4_START_ADDR                  => 23040,
			SECTOR4_END_ADDR                    => 58879,
			SECTOR5_START_ADDR                  => 0,
			SECTOR5_END_ADDR                    => 0,
			MIN_VALID_ADDR                      => 0,
			MAX_VALID_ADDR                      => 58879,
			MIN_UFM_VALID_ADDR                  => 0,
			MAX_UFM_VALID_ADDR                  => 8191,
			SECTOR1_MAP                         => 1,
			SECTOR2_MAP                         => 2,
			SECTOR3_MAP                         => 4,
			SECTOR4_MAP                         => 5,
			SECTOR5_MAP                         => 0,
			ADDR_RANGE1_END_ADDR                => 8191,
			ADDR_RANGE1_OFFSET                  => 512,
			ADDR_RANGE2_OFFSET                  => 21504,
			AVMM_DATA_ADDR_WIDTH                => 16,
			AVMM_DATA_DATA_WIDTH                => 32,
			AVMM_DATA_BURSTCOUNT_WIDTH          => 4,
			SECTOR_READ_PROTECTION_MODE         => 16,
			FLASH_SEQ_READ_DATA_COUNT           => 2,
			FLASH_ADDR_ALIGNMENT_BITS           => 1,
			FLASH_READ_CYCLE_MAX_INDEX          => 4,
			FLASH_RESET_CYCLE_MAX_INDEX         => 28,
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  => 135,
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX => 39516766,
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX => 34436,
			PARALLEL_MODE                       => true,
			READ_AND_WRITE_MODE                 => true,
			WRAPPING_BURST_MODE                 => false,
			IS_DUAL_BOOT                        => "False",
			IS_ERAM_SKIP                        => "True",
			IS_COMPRESSED_IMAGE                 => "False"
		)
		port map (
			clock                   => altpll_0_c0_clk,                                     --    clk.clk
			reset_n                 => rst_controller_reset_out_reset_ports_inv,            -- nreset.reset_n
			avmm_data_addr          => mm_interconnect_0_onchip_flash_0_data_address,       --   data.address
			avmm_data_read          => mm_interconnect_0_onchip_flash_0_data_read,          --       .read
			avmm_data_writedata     => mm_interconnect_0_onchip_flash_0_data_writedata,     --       .writedata
			avmm_data_write         => mm_interconnect_0_onchip_flash_0_data_write,         --       .write
			avmm_data_readdata      => mm_interconnect_0_onchip_flash_0_data_readdata,      --       .readdata
			avmm_data_waitrequest   => mm_interconnect_0_onchip_flash_0_data_waitrequest,   --       .waitrequest
			avmm_data_readdatavalid => mm_interconnect_0_onchip_flash_0_data_readdatavalid, --       .readdatavalid
			avmm_data_burstcount    => mm_interconnect_0_onchip_flash_0_data_burstcount,    --       .burstcount
			avmm_csr_addr           => mm_interconnect_0_onchip_flash_0_csr_address(0),     --    csr.address
			avmm_csr_read           => mm_interconnect_0_onchip_flash_0_csr_read,           --       .read
			avmm_csr_writedata      => mm_interconnect_0_onchip_flash_0_csr_writedata,      --       .writedata
			avmm_csr_write          => mm_interconnect_0_onchip_flash_0_csr_write,          --       .write
			avmm_csr_readdata       => mm_interconnect_0_onchip_flash_0_csr_readdata        --       .readdata
		);

	onchip_memory2_0 : component wasca_onchip_memory2_0
		port map (
			clk        => altpll_0_c0_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                --       .reset_req
		);

	onchip_memory2_1 : component wasca_onchip_memory2_1
		port map (
			clk        => altpll_0_c0_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_1_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_1_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_1_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_1_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_1_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_1_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_1_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                --       .reset_req
		);

	performance_counter_0 : component wasca_performance_counter_0
		port map (
			clk           => altpll_0_c0_clk,                                                     --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                            --         reset.reset_n
			address       => mm_interconnect_0_performance_counter_0_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_performance_counter_0_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_performance_counter_0_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_performance_counter_0_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_performance_counter_0_control_slave_writedata      --              .writedata
		);

	switches : component wasca_switches
		port map (
			clk      => altpll_0_c0_clk,                          --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switches_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_switches_s1_readdata,   --                    .readdata
			in_port  => switches_conn_export                      -- external_connection.export
		);

	uart_0 : component wasca_uart_0
		port map (
			clk           => altpll_0_c0_clk,                             --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_0_uart_0_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_0_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_0_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_0_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_0_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_0_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_0_s1_readdata,        --                    .readdata
			dataavailable => open,                                        --                    .dataavailable
			readyfordata  => open,                                        --                    .readyfordata
			rxd           => uart_0_external_connection_rxd,              -- external_connection.export
			txd           => uart_0_external_connection_txd,              --                    .export
			irq           => irq_mapper_receiver0_irq                     --                 irq.irq
		);

	mm_interconnect_0 : component wasca_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                            => altpll_0_c0_clk,                                                     --                                          altpll_0_c0.clk
			clk_0_clk_clk                                              => clk_clk,                                                             --                                            clk_0_clk.clk
			abus_slave_0_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                                      --             abus_slave_0_reset_reset_bridge_in_reset.reset
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                  -- altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			abus_slave_0_avalon_master_address                         => abus_slave_0_avalon_master_address,                                  --                           abus_slave_0_avalon_master.address
			abus_slave_0_avalon_master_waitrequest                     => abus_slave_0_avalon_master_waitrequest,                              --                                                     .waitrequest
			abus_slave_0_avalon_master_burstcount(0)                   => abus_slave_0_avalon_master_burstcount,                               --                                                     .burstcount
			abus_slave_0_avalon_master_read                            => abus_slave_0_avalon_master_read,                                     --                                                     .read
			abus_slave_0_avalon_master_readdata                        => abus_slave_0_avalon_master_readdata,                                 --                                                     .readdata
			abus_slave_0_avalon_master_readdatavalid                   => abus_slave_0_avalon_master_readdatavalid,                            --                                                     .readdatavalid
			abus_slave_0_avalon_master_write                           => abus_slave_0_avalon_master_write,                                    --                                                     .write
			abus_slave_0_avalon_master_writedata                       => abus_slave_0_avalon_master_writedata,                                --                                                     .writedata
			nios2_gen2_0_data_master_address                           => nios2_gen2_0_data_master_address,                                    --                             nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                                --                                                     .waitrequest
			nios2_gen2_0_data_master_byteenable                        => nios2_gen2_0_data_master_byteenable,                                 --                                                     .byteenable
			nios2_gen2_0_data_master_read                              => nios2_gen2_0_data_master_read,                                       --                                                     .read
			nios2_gen2_0_data_master_readdata                          => nios2_gen2_0_data_master_readdata,                                   --                                                     .readdata
			nios2_gen2_0_data_master_write                             => nios2_gen2_0_data_master_write,                                      --                                                     .write
			nios2_gen2_0_data_master_writedata                         => nios2_gen2_0_data_master_writedata,                                  --                                                     .writedata
			nios2_gen2_0_data_master_debugaccess                       => nios2_gen2_0_data_master_debugaccess,                                --                                                     .debugaccess
			nios2_gen2_0_instruction_master_address                    => nios2_gen2_0_instruction_master_address,                             --                      nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                => nios2_gen2_0_instruction_master_waitrequest,                         --                                                     .waitrequest
			nios2_gen2_0_instruction_master_read                       => nios2_gen2_0_instruction_master_read,                                --                                                     .read
			nios2_gen2_0_instruction_master_readdata                   => nios2_gen2_0_instruction_master_readdata,                            --                                                     .readdata
			abus_demux_0_avalon_nios_address                           => mm_interconnect_0_abus_demux_0_avalon_nios_address,                  --                             abus_demux_0_avalon_nios.address
			abus_demux_0_avalon_nios_write                             => mm_interconnect_0_abus_demux_0_avalon_nios_write,                    --                                                     .write
			abus_demux_0_avalon_nios_read                              => mm_interconnect_0_abus_demux_0_avalon_nios_read,                     --                                                     .read
			abus_demux_0_avalon_nios_readdata                          => mm_interconnect_0_abus_demux_0_avalon_nios_readdata,                 --                                                     .readdata
			abus_demux_0_avalon_nios_writedata                         => mm_interconnect_0_abus_demux_0_avalon_nios_writedata,                --                                                     .writedata
			abus_demux_0_avalon_nios_burstcount                        => mm_interconnect_0_abus_demux_0_avalon_nios_burstcount,               --                                                     .burstcount
			abus_demux_0_avalon_nios_readdatavalid                     => mm_interconnect_0_abus_demux_0_avalon_nios_readdatavalid,            --                                                     .readdatavalid
			abus_demux_0_avalon_nios_waitrequest                       => mm_interconnect_0_abus_demux_0_avalon_nios_waitrequest,              --                                                     .waitrequest
			abus_slave_0_avalon_nios_address                           => mm_interconnect_0_abus_slave_0_avalon_nios_address,                  --                             abus_slave_0_avalon_nios.address
			abus_slave_0_avalon_nios_write                             => mm_interconnect_0_abus_slave_0_avalon_nios_write,                    --                                                     .write
			abus_slave_0_avalon_nios_read                              => mm_interconnect_0_abus_slave_0_avalon_nios_read,                     --                                                     .read
			abus_slave_0_avalon_nios_readdata                          => mm_interconnect_0_abus_slave_0_avalon_nios_readdata,                 --                                                     .readdata
			abus_slave_0_avalon_nios_writedata                         => mm_interconnect_0_abus_slave_0_avalon_nios_writedata,                --                                                     .writedata
			abus_slave_0_avalon_nios_burstcount                        => mm_interconnect_0_abus_slave_0_avalon_nios_burstcount,               --                                                     .burstcount
			abus_slave_0_avalon_nios_readdatavalid                     => mm_interconnect_0_abus_slave_0_avalon_nios_readdatavalid,            --                                                     .readdatavalid
			abus_slave_0_avalon_nios_waitrequest                       => mm_interconnect_0_abus_slave_0_avalon_nios_waitrequest,              --                                                     .waitrequest
			altpll_0_pll_slave_address                                 => mm_interconnect_0_altpll_0_pll_slave_address,                        --                                   altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                   => mm_interconnect_0_altpll_0_pll_slave_write,                          --                                                     .write
			altpll_0_pll_slave_read                                    => mm_interconnect_0_altpll_0_pll_slave_read,                           --                                                     .read
			altpll_0_pll_slave_readdata                                => mm_interconnect_0_altpll_0_pll_slave_readdata,                       --                                                     .readdata
			altpll_0_pll_slave_writedata                               => mm_interconnect_0_altpll_0_pll_slave_writedata,                      --                                                     .writedata
			external_sdram_controller_s1_address                       => mm_interconnect_0_external_sdram_controller_s1_address,              --                         external_sdram_controller_s1.address
			external_sdram_controller_s1_write                         => mm_interconnect_0_external_sdram_controller_s1_write,                --                                                     .write
			external_sdram_controller_s1_read                          => mm_interconnect_0_external_sdram_controller_s1_read,                 --                                                     .read
			external_sdram_controller_s1_readdata                      => mm_interconnect_0_external_sdram_controller_s1_readdata,             --                                                     .readdata
			external_sdram_controller_s1_writedata                     => mm_interconnect_0_external_sdram_controller_s1_writedata,            --                                                     .writedata
			external_sdram_controller_s1_byteenable                    => mm_interconnect_0_external_sdram_controller_s1_byteenable,           --                                                     .byteenable
			external_sdram_controller_s1_readdatavalid                 => mm_interconnect_0_external_sdram_controller_s1_readdatavalid,        --                                                     .readdatavalid
			external_sdram_controller_s1_waitrequest                   => mm_interconnect_0_external_sdram_controller_s1_waitrequest,          --                                                     .waitrequest
			external_sdram_controller_s1_chipselect                    => mm_interconnect_0_external_sdram_controller_s1_chipselect,           --                                                     .chipselect
			leds_s1_address                                            => mm_interconnect_0_leds_s1_address,                                   --                                              leds_s1.address
			leds_s1_write                                              => mm_interconnect_0_leds_s1_write,                                     --                                                     .write
			leds_s1_readdata                                           => mm_interconnect_0_leds_s1_readdata,                                  --                                                     .readdata
			leds_s1_writedata                                          => mm_interconnect_0_leds_s1_writedata,                                 --                                                     .writedata
			leds_s1_chipselect                                         => mm_interconnect_0_leds_s1_chipselect,                                --                                                     .chipselect
			nios2_gen2_0_debug_mem_slave_address                       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,              --                         nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                --                                                     .write
			nios2_gen2_0_debug_mem_slave_read                          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                 --                                                     .read
			nios2_gen2_0_debug_mem_slave_readdata                      => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,             --                                                     .readdata
			nios2_gen2_0_debug_mem_slave_writedata                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,            --                                                     .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,           --                                                     .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,          --                                                     .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,          --                                                     .debugaccess
			onchip_flash_0_csr_address                                 => mm_interconnect_0_onchip_flash_0_csr_address,                        --                                   onchip_flash_0_csr.address
			onchip_flash_0_csr_write                                   => mm_interconnect_0_onchip_flash_0_csr_write,                          --                                                     .write
			onchip_flash_0_csr_read                                    => mm_interconnect_0_onchip_flash_0_csr_read,                           --                                                     .read
			onchip_flash_0_csr_readdata                                => mm_interconnect_0_onchip_flash_0_csr_readdata,                       --                                                     .readdata
			onchip_flash_0_csr_writedata                               => mm_interconnect_0_onchip_flash_0_csr_writedata,                      --                                                     .writedata
			onchip_flash_0_data_address                                => mm_interconnect_0_onchip_flash_0_data_address,                       --                                  onchip_flash_0_data.address
			onchip_flash_0_data_write                                  => mm_interconnect_0_onchip_flash_0_data_write,                         --                                                     .write
			onchip_flash_0_data_read                                   => mm_interconnect_0_onchip_flash_0_data_read,                          --                                                     .read
			onchip_flash_0_data_readdata                               => mm_interconnect_0_onchip_flash_0_data_readdata,                      --                                                     .readdata
			onchip_flash_0_data_writedata                              => mm_interconnect_0_onchip_flash_0_data_writedata,                     --                                                     .writedata
			onchip_flash_0_data_burstcount                             => mm_interconnect_0_onchip_flash_0_data_burstcount,                    --                                                     .burstcount
			onchip_flash_0_data_readdatavalid                          => mm_interconnect_0_onchip_flash_0_data_readdatavalid,                 --                                                     .readdatavalid
			onchip_flash_0_data_waitrequest                            => mm_interconnect_0_onchip_flash_0_data_waitrequest,                   --                                                     .waitrequest
			onchip_memory2_0_s1_address                                => mm_interconnect_0_onchip_memory2_0_s1_address,                       --                                  onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                  => mm_interconnect_0_onchip_memory2_0_s1_write,                         --                                                     .write
			onchip_memory2_0_s1_readdata                               => mm_interconnect_0_onchip_memory2_0_s1_readdata,                      --                                                     .readdata
			onchip_memory2_0_s1_writedata                              => mm_interconnect_0_onchip_memory2_0_s1_writedata,                     --                                                     .writedata
			onchip_memory2_0_s1_byteenable                             => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                    --                                                     .byteenable
			onchip_memory2_0_s1_chipselect                             => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                    --                                                     .chipselect
			onchip_memory2_0_s1_clken                                  => mm_interconnect_0_onchip_memory2_0_s1_clken,                         --                                                     .clken
			onchip_memory2_1_s1_address                                => mm_interconnect_0_onchip_memory2_1_s1_address,                       --                                  onchip_memory2_1_s1.address
			onchip_memory2_1_s1_write                                  => mm_interconnect_0_onchip_memory2_1_s1_write,                         --                                                     .write
			onchip_memory2_1_s1_readdata                               => mm_interconnect_0_onchip_memory2_1_s1_readdata,                      --                                                     .readdata
			onchip_memory2_1_s1_writedata                              => mm_interconnect_0_onchip_memory2_1_s1_writedata,                     --                                                     .writedata
			onchip_memory2_1_s1_byteenable                             => mm_interconnect_0_onchip_memory2_1_s1_byteenable,                    --                                                     .byteenable
			onchip_memory2_1_s1_chipselect                             => mm_interconnect_0_onchip_memory2_1_s1_chipselect,                    --                                                     .chipselect
			onchip_memory2_1_s1_clken                                  => mm_interconnect_0_onchip_memory2_1_s1_clken,                         --                                                     .clken
			performance_counter_0_control_slave_address                => mm_interconnect_0_performance_counter_0_control_slave_address,       --                  performance_counter_0_control_slave.address
			performance_counter_0_control_slave_write                  => mm_interconnect_0_performance_counter_0_control_slave_write,         --                                                     .write
			performance_counter_0_control_slave_readdata               => mm_interconnect_0_performance_counter_0_control_slave_readdata,      --                                                     .readdata
			performance_counter_0_control_slave_writedata              => mm_interconnect_0_performance_counter_0_control_slave_writedata,     --                                                     .writedata
			performance_counter_0_control_slave_begintransfer          => mm_interconnect_0_performance_counter_0_control_slave_begintransfer, --                                                     .begintransfer
			switches_s1_address                                        => mm_interconnect_0_switches_s1_address,                               --                                          switches_s1.address
			switches_s1_readdata                                       => mm_interconnect_0_switches_s1_readdata,                              --                                                     .readdata
			uart_0_s1_address                                          => mm_interconnect_0_uart_0_s1_address,                                 --                                            uart_0_s1.address
			uart_0_s1_write                                            => mm_interconnect_0_uart_0_s1_write,                                   --                                                     .write
			uart_0_s1_read                                             => mm_interconnect_0_uart_0_s1_read,                                    --                                                     .read
			uart_0_s1_readdata                                         => mm_interconnect_0_uart_0_s1_readdata,                                --                                                     .readdata
			uart_0_s1_writedata                                        => mm_interconnect_0_uart_0_s1_writedata,                               --                                                     .writedata
			uart_0_s1_begintransfer                                    => mm_interconnect_0_uart_0_s1_begintransfer,                           --                                                     .begintransfer
			uart_0_s1_chipselect                                       => mm_interconnect_0_uart_0_s1_chipselect                               --                                                     .chipselect
		);

	irq_mapper : component wasca_irq_mapper
		port map (
			clk           => altpll_0_c0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component wasca_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			clk            => altpll_0_c0_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component wasca_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component wasca_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "both",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_gen2_0_debug_reset_request_reset, -- reset_in0.reset
			clk            => altpll_0_c0_clk,                        --       clk.clk
			reset_out      => open,                                   -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_external_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_external_sdram_controller_s1_read;

	mm_interconnect_0_external_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_external_sdram_controller_s1_byteenable;

	mm_interconnect_0_external_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_external_sdram_controller_s1_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_uart_0_s1_read_ports_inv <= not mm_interconnect_0_uart_0_s1_read;

	mm_interconnect_0_uart_0_s1_write_ports_inv <= not mm_interconnect_0_uart_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	clock_116_mhz_clk <= altpll_0_c0_clk;

end architecture rtl; -- of wasca
