// wasca.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module wasca (
		input  wire [9:0]  abus_avalon_sdram_bridge_0_abus_address,           //  abus_avalon_sdram_bridge_0_abus.address
		input  wire        abus_avalon_sdram_bridge_0_abus_read,              //                                 .read
		output wire        abus_avalon_sdram_bridge_0_abus_waitrequest,       //                                 .waitrequest
		inout  wire [15:0] abus_avalon_sdram_bridge_0_abus_addressdata,       //                                 .addressdata
		input  wire [2:0]  abus_avalon_sdram_bridge_0_abus_chipselect,        //                                 .chipselect
		output wire        abus_avalon_sdram_bridge_0_abus_direction,         //                                 .direction
		output wire        abus_avalon_sdram_bridge_0_abus_disable_out,       //                                 .disable_out
		output wire        abus_avalon_sdram_bridge_0_abus_interrupt,         //                                 .interrupt
		output wire [1:0]  abus_avalon_sdram_bridge_0_abus_muxing,            //                                 .muxing
		input  wire [1:0]  abus_avalon_sdram_bridge_0_abus_writebyteenable_n, //                                 .writebyteenable_n
		input  wire        abus_avalon_sdram_bridge_0_abus_reset,             //                                 .reset
		output wire [12:0] abus_avalon_sdram_bridge_0_sdram_addr,             // abus_avalon_sdram_bridge_0_sdram.addr
		output wire [1:0]  abus_avalon_sdram_bridge_0_sdram_ba,               //                                 .ba
		output wire        abus_avalon_sdram_bridge_0_sdram_cas_n,            //                                 .cas_n
		output wire        abus_avalon_sdram_bridge_0_sdram_cke,              //                                 .cke
		output wire        abus_avalon_sdram_bridge_0_sdram_cs_n,             //                                 .cs_n
		inout  wire [15:0] abus_avalon_sdram_bridge_0_sdram_dq,               //                                 .dq
		output wire [1:0]  abus_avalon_sdram_bridge_0_sdram_dqm,              //                                 .dqm
		output wire        abus_avalon_sdram_bridge_0_sdram_ras_n,            //                                 .ras_n
		output wire        abus_avalon_sdram_bridge_0_sdram_we_n,             //                                 .we_n
		output wire        abus_avalon_sdram_bridge_0_sdram_clk,              //                                 .clk
		input  wire        altpll_1_areset_conduit_export,                    //          altpll_1_areset_conduit.export
		output wire        altpll_1_locked_conduit_export,                    //          altpll_1_locked_conduit.export
		output wire        altpll_1_phasedone_conduit_export,                 //       altpll_1_phasedone_conduit.export
		output wire        buffered_spi_mosi,                                 //                     buffered_spi.mosi
		output wire        buffered_spi_clk,                                  //                                 .clk
		input  wire        buffered_spi_miso,                                 //                                 .miso
		output wire        buffered_spi_cs,                                   //                                 .cs
		input  wire        clk_clk,                                           //                              clk.clk
		output wire        clock_116_mhz_clk,                                 //                    clock_116_mhz.clk
		output wire [4:0]  extra_leds_conn_export,                            //                  extra_leds_conn.export
		output wire [6:0]  hex0_conn_export,                                  //                        hex0_conn.export
		output wire [6:0]  hex1_conn_export,                                  //                        hex1_conn.export
		output wire [6:0]  hex2_conn_export,                                  //                        hex2_conn.export
		output wire [6:0]  hex3_conn_export,                                  //                        hex3_conn.export
		output wire [6:0]  hex4_conn_export,                                  //                        hex4_conn.export
		output wire [6:0]  hex5_conn_export,                                  //                        hex5_conn.export
		output wire [5:0]  hexdot_conn_export,                                //                      hexdot_conn.export
		output wire [3:0]  leds_conn_export,                                  //                        leds_conn.export
		input  wire        reset_reset_n,                                     //                            reset.reset_n
		input  wire        reset_controller_0_reset_in1_reset,                //     reset_controller_0_reset_in1.reset
		input  wire        spi_sync_conn_export,                              //                    spi_sync_conn.export
		input  wire [7:0]  switches_conn_export,                              //                    switches_conn.export
		input  wire        uart_0_external_connection_rxd,                    //       uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd                     //                                 .txd
	);

	wire         nios2_gen2_0_debug_reset_request_reset;                                  // nios2_gen2_0:debug_reset_request -> [buffered_spi_0:reset, extra_leds:reset_n, hex0:reset_n, hex1:reset_n, hex2:reset_n, hex3:reset_n, hex4:reset_n, hex5:reset_n, hexdot:reset_n, leds:reset_n, mm_interconnect_0:buffered_spi_0_reset_reset_bridge_in_reset_reset, performance_counter_0:reset_n, reset_controller_0:reset_in0, spi_sync:reset_n, switches:reset_n]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                       // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                    // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                    // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                                        // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                     // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                           // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                          // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                      // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                             // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [24:0] nios2_gen2_0_instruction_master_address;                                 // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                    // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [15:0] mm_interconnect_0_buffered_spi_0_avalon_readdata;                        // buffered_spi_0:avalon_readdata -> mm_interconnect_0:buffered_spi_0_avalon_readdata
	wire         mm_interconnect_0_buffered_spi_0_avalon_waitrequest;                     // buffered_spi_0:avalon_waitrequest -> mm_interconnect_0:buffered_spi_0_avalon_waitrequest
	wire  [13:0] mm_interconnect_0_buffered_spi_0_avalon_address;                         // mm_interconnect_0:buffered_spi_0_avalon_address -> buffered_spi_0:avalon_address
	wire         mm_interconnect_0_buffered_spi_0_avalon_read;                            // mm_interconnect_0:buffered_spi_0_avalon_read -> buffered_spi_0:avalon_read
	wire         mm_interconnect_0_buffered_spi_0_avalon_readdatavalid;                   // buffered_spi_0:avalon_readdatavalid -> mm_interconnect_0:buffered_spi_0_avalon_readdatavalid
	wire         mm_interconnect_0_buffered_spi_0_avalon_write;                           // mm_interconnect_0:buffered_spi_0_avalon_write -> buffered_spi_0:avalon_write
	wire  [15:0] mm_interconnect_0_buffered_spi_0_avalon_writedata;                       // mm_interconnect_0:buffered_spi_0_avalon_writedata -> buffered_spi_0:avalon_writedata
	wire  [15:0] mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_readdata;       // abus_avalon_sdram_bridge_0:avalon_regs_readdata -> mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_regs_readdata
	wire         mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_waitrequest;    // abus_avalon_sdram_bridge_0:avalon_regs_waitrequest -> mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_regs_waitrequest
	wire   [7:0] mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_address;        // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_regs_address -> abus_avalon_sdram_bridge_0:avalon_regs_address
	wire         mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_read;           // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_regs_read -> abus_avalon_sdram_bridge_0:avalon_regs_read
	wire         mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_readdatavalid;  // abus_avalon_sdram_bridge_0:avalon_regs_readdatavalid -> mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_regs_readdatavalid
	wire         mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_write;          // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_regs_write -> abus_avalon_sdram_bridge_0:avalon_regs_write
	wire  [15:0] mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_writedata;      // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_regs_writedata -> abus_avalon_sdram_bridge_0:avalon_regs_writedata
	wire  [15:0] mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_readdata;      // abus_avalon_sdram_bridge_0:avalon_sdram_readdata -> mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_sdram_readdata
	wire         mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_waitrequest;   // abus_avalon_sdram_bridge_0:avalon_sdram_waitrequest -> mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_sdram_waitrequest
	wire  [24:0] mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_address;       // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_sdram_address -> abus_avalon_sdram_bridge_0:avalon_sdram_address
	wire         mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_read;          // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_sdram_read -> abus_avalon_sdram_bridge_0:avalon_sdram_read
	wire   [1:0] mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_byteenable;    // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_sdram_byteenable -> abus_avalon_sdram_bridge_0:avalon_sdram_byteenable
	wire         mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_readdatavalid; // abus_avalon_sdram_bridge_0:avalon_sdram_readdatavalid -> mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_sdram_readdatavalid
	wire         mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_write;         // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_sdram_write -> abus_avalon_sdram_bridge_0:avalon_sdram_write
	wire  [15:0] mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_writedata;     // mm_interconnect_0:abus_avalon_sdram_bridge_0_avalon_sdram_writedata -> abus_avalon_sdram_bridge_0:avalon_sdram_writedata
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_readdata;          // performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	wire   [2:0] mm_interconnect_0_performance_counter_0_control_slave_address;           // mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	wire         mm_interconnect_0_performance_counter_0_control_slave_begintransfer;     // mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	wire         mm_interconnect_0_performance_counter_0_control_slave_write;             // mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_writedata;         // mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_readdata;                           // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	wire   [0:0] mm_interconnect_0_onchip_flash_0_csr_address;                            // mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_0_onchip_flash_0_csr_read;                               // mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire         mm_interconnect_0_onchip_flash_0_csr_write;                              // mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_writedata;                          // mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;                          // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;                       // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire  [18:0] mm_interconnect_0_onchip_flash_0_data_address;                           // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_read;                              // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;                     // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_onchip_flash_0_data_write;                             // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;                         // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;                        // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                 // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;              // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;               // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_1_pll_slave_readdata;                           // altpll_1:readdata -> mm_interconnect_0:altpll_1_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_1_pll_slave_address;                            // mm_interconnect_0:altpll_1_pll_slave_address -> altpll_1:address
	wire         mm_interconnect_0_altpll_1_pll_slave_read;                               // mm_interconnect_0:altpll_1_pll_slave_read -> altpll_1:read
	wire         mm_interconnect_0_altpll_1_pll_slave_write;                              // mm_interconnect_0:altpll_1_pll_slave_write -> altpll_1:write
	wire  [31:0] mm_interconnect_0_altpll_1_pll_slave_writedata;                          // mm_interconnect_0:altpll_1_pll_slave_writedata -> altpll_1:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                        // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                          // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;                           // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                        // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                             // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                         // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                             // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_uart_0_s1_chipselect;                                  // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                                    // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                     // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                        // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                               // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                       // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                                   // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                                  // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                                   // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                    // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                      // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                       // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                         // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                     // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_extra_leds_s1_chipselect;                              // mm_interconnect_0:extra_leds_s1_chipselect -> extra_leds:chipselect
	wire  [31:0] mm_interconnect_0_extra_leds_s1_readdata;                                // extra_leds:readdata -> mm_interconnect_0:extra_leds_s1_readdata
	wire   [1:0] mm_interconnect_0_extra_leds_s1_address;                                 // mm_interconnect_0:extra_leds_s1_address -> extra_leds:address
	wire         mm_interconnect_0_extra_leds_s1_write;                                   // mm_interconnect_0:extra_leds_s1_write -> extra_leds:write_n
	wire  [31:0] mm_interconnect_0_extra_leds_s1_writedata;                               // mm_interconnect_0:extra_leds_s1_writedata -> extra_leds:writedata
	wire         mm_interconnect_0_hex0_s1_chipselect;                                    // mm_interconnect_0:hex0_s1_chipselect -> hex0:chipselect
	wire  [31:0] mm_interconnect_0_hex0_s1_readdata;                                      // hex0:readdata -> mm_interconnect_0:hex0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_s1_address;                                       // mm_interconnect_0:hex0_s1_address -> hex0:address
	wire         mm_interconnect_0_hex0_s1_write;                                         // mm_interconnect_0:hex0_s1_write -> hex0:write_n
	wire  [31:0] mm_interconnect_0_hex0_s1_writedata;                                     // mm_interconnect_0:hex0_s1_writedata -> hex0:writedata
	wire         mm_interconnect_0_hex1_s1_chipselect;                                    // mm_interconnect_0:hex1_s1_chipselect -> hex1:chipselect
	wire  [31:0] mm_interconnect_0_hex1_s1_readdata;                                      // hex1:readdata -> mm_interconnect_0:hex1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex1_s1_address;                                       // mm_interconnect_0:hex1_s1_address -> hex1:address
	wire         mm_interconnect_0_hex1_s1_write;                                         // mm_interconnect_0:hex1_s1_write -> hex1:write_n
	wire  [31:0] mm_interconnect_0_hex1_s1_writedata;                                     // mm_interconnect_0:hex1_s1_writedata -> hex1:writedata
	wire         mm_interconnect_0_hex2_s1_chipselect;                                    // mm_interconnect_0:hex2_s1_chipselect -> hex2:chipselect
	wire  [31:0] mm_interconnect_0_hex2_s1_readdata;                                      // hex2:readdata -> mm_interconnect_0:hex2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex2_s1_address;                                       // mm_interconnect_0:hex2_s1_address -> hex2:address
	wire         mm_interconnect_0_hex2_s1_write;                                         // mm_interconnect_0:hex2_s1_write -> hex2:write_n
	wire  [31:0] mm_interconnect_0_hex2_s1_writedata;                                     // mm_interconnect_0:hex2_s1_writedata -> hex2:writedata
	wire         mm_interconnect_0_hex3_s1_chipselect;                                    // mm_interconnect_0:hex3_s1_chipselect -> hex3:chipselect
	wire  [31:0] mm_interconnect_0_hex3_s1_readdata;                                      // hex3:readdata -> mm_interconnect_0:hex3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_s1_address;                                       // mm_interconnect_0:hex3_s1_address -> hex3:address
	wire         mm_interconnect_0_hex3_s1_write;                                         // mm_interconnect_0:hex3_s1_write -> hex3:write_n
	wire  [31:0] mm_interconnect_0_hex3_s1_writedata;                                     // mm_interconnect_0:hex3_s1_writedata -> hex3:writedata
	wire         mm_interconnect_0_hex5_s1_chipselect;                                    // mm_interconnect_0:hex5_s1_chipselect -> hex5:chipselect
	wire  [31:0] mm_interconnect_0_hex5_s1_readdata;                                      // hex5:readdata -> mm_interconnect_0:hex5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_s1_address;                                       // mm_interconnect_0:hex5_s1_address -> hex5:address
	wire         mm_interconnect_0_hex5_s1_write;                                         // mm_interconnect_0:hex5_s1_write -> hex5:write_n
	wire  [31:0] mm_interconnect_0_hex5_s1_writedata;                                     // mm_interconnect_0:hex5_s1_writedata -> hex5:writedata
	wire         mm_interconnect_0_hex4_s1_chipselect;                                    // mm_interconnect_0:hex4_s1_chipselect -> hex4:chipselect
	wire  [31:0] mm_interconnect_0_hex4_s1_readdata;                                      // hex4:readdata -> mm_interconnect_0:hex4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_s1_address;                                       // mm_interconnect_0:hex4_s1_address -> hex4:address
	wire         mm_interconnect_0_hex4_s1_write;                                         // mm_interconnect_0:hex4_s1_write -> hex4:write_n
	wire  [31:0] mm_interconnect_0_hex4_s1_writedata;                                     // mm_interconnect_0:hex4_s1_writedata -> hex4:writedata
	wire         mm_interconnect_0_hexdot_s1_chipselect;                                  // mm_interconnect_0:hexdot_s1_chipselect -> hexdot:chipselect
	wire  [31:0] mm_interconnect_0_hexdot_s1_readdata;                                    // hexdot:readdata -> mm_interconnect_0:hexdot_s1_readdata
	wire   [1:0] mm_interconnect_0_hexdot_s1_address;                                     // mm_interconnect_0:hexdot_s1_address -> hexdot:address
	wire         mm_interconnect_0_hexdot_s1_write;                                       // mm_interconnect_0:hexdot_s1_write -> hexdot:write_n
	wire  [31:0] mm_interconnect_0_hexdot_s1_writedata;                                   // mm_interconnect_0:hexdot_s1_writedata -> hexdot:writedata
	wire  [31:0] mm_interconnect_0_spi_sync_s1_readdata;                                  // spi_sync:readdata -> mm_interconnect_0:spi_sync_s1_readdata
	wire   [1:0] mm_interconnect_0_spi_sync_s1_address;                                   // mm_interconnect_0:spi_sync_s1_address -> spi_sync:address
	wire         irq_mapper_receiver0_irq;                                                // uart_0:irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                    // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [abus_avalon_sdram_bridge_0:reset, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_flash_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         reset_controller_0_reset_out_reset;                                      // reset_controller_0:reset_out -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [altpll_1:reset, mm_interconnect_0:altpll_1_inclk_interface_reset_reset_bridge_in_reset_reset]

	abus_avalon_sdram_bridge abus_avalon_sdram_bridge_0 (
		.abus_address               (abus_avalon_sdram_bridge_0_abus_address),                                 //         abus.address
		.abus_read                  (abus_avalon_sdram_bridge_0_abus_read),                                    //             .read
		.abus_waitrequest           (abus_avalon_sdram_bridge_0_abus_waitrequest),                             //             .waitrequest
		.abus_addressdata           (abus_avalon_sdram_bridge_0_abus_addressdata),                             //             .addressdata
		.abus_chipselect            (abus_avalon_sdram_bridge_0_abus_chipselect),                              //             .chipselect
		.abus_direction             (abus_avalon_sdram_bridge_0_abus_direction),                               //             .direction
		.abus_disable_out           (abus_avalon_sdram_bridge_0_abus_disable_out),                             //             .disable_out
		.abus_interrupt             (abus_avalon_sdram_bridge_0_abus_interrupt),                               //             .interrupt
		.abus_muxing                (abus_avalon_sdram_bridge_0_abus_muxing),                                  //             .muxing
		.abus_write                 (abus_avalon_sdram_bridge_0_abus_writebyteenable_n),                       //             .writebyteenable_n
		.saturn_reset               (abus_avalon_sdram_bridge_0_abus_reset),                                   //             .reset
		.avalon_sdram_read          (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_read),          // avalon_sdram.read
		.avalon_sdram_write         (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_write),         //             .write
		.avalon_sdram_waitrequest   (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_waitrequest),   //             .waitrequest
		.avalon_sdram_address       (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_address),       //             .address
		.avalon_sdram_writedata     (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_writedata),     //             .writedata
		.avalon_sdram_readdata      (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_readdata),      //             .readdata
		.avalon_sdram_readdatavalid (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_readdatavalid), //             .readdatavalid
		.avalon_sdram_byteenable    (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_byteenable),    //             .byteenable
		.avalon_regs_read           (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_read),           //  avalon_regs.read
		.avalon_regs_write          (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_write),          //             .write
		.avalon_regs_waitrequest    (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_waitrequest),    //             .waitrequest
		.avalon_regs_address        (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_address),        //             .address
		.avalon_regs_writedata      (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_writedata),      //             .writedata
		.avalon_regs_readdata       (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_readdata),       //             .readdata
		.avalon_regs_readdatavalid  (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_readdatavalid),  //             .readdatavalid
		.reset                      (rst_controller_reset_out_reset),                                          //        reset.reset
		.clock                      (clock_116_mhz_clk),                                                       //        clock.clk
		.sdram_addr                 (abus_avalon_sdram_bridge_0_sdram_addr),                                   //        sdram.addr
		.sdram_ba                   (abus_avalon_sdram_bridge_0_sdram_ba),                                     //             .ba
		.sdram_cas_n                (abus_avalon_sdram_bridge_0_sdram_cas_n),                                  //             .cas_n
		.sdram_cke                  (abus_avalon_sdram_bridge_0_sdram_cke),                                    //             .cke
		.sdram_cs_n                 (abus_avalon_sdram_bridge_0_sdram_cs_n),                                   //             .cs_n
		.sdram_dq                   (abus_avalon_sdram_bridge_0_sdram_dq),                                     //             .dq
		.sdram_dqm                  (abus_avalon_sdram_bridge_0_sdram_dqm),                                    //             .dqm
		.sdram_ras_n                (abus_avalon_sdram_bridge_0_sdram_ras_n),                                  //             .ras_n
		.sdram_we_n                 (abus_avalon_sdram_bridge_0_sdram_we_n),                                   //             .we_n
		.sdram_clk                  (abus_avalon_sdram_bridge_0_sdram_clk)                                     //             .clk
	);

	wasca_altpll_1 altpll_1 (
		.clk       (clk_clk),                                        //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_1_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_1_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_1_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_1_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_1_pll_slave_writedata), //                      .writedata
		.c0        (clock_116_mhz_clk),                              //                    c0.clk
		.areset    (altpll_1_areset_conduit_export),                 //        areset_conduit.export
		.locked    (altpll_1_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_1_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	buffered_spi buffered_spi_0 (
		.reset                (nios2_gen2_0_debug_reset_request_reset),                //       reset.reset
		.avalon_read          (mm_interconnect_0_buffered_spi_0_avalon_read),          //      avalon.read
		.avalon_write         (mm_interconnect_0_buffered_spi_0_avalon_write),         //            .write
		.avalon_address       (mm_interconnect_0_buffered_spi_0_avalon_address),       //            .address
		.avalon_waitrequest   (mm_interconnect_0_buffered_spi_0_avalon_waitrequest),   //            .waitrequest
		.avalon_writedata     (mm_interconnect_0_buffered_spi_0_avalon_writedata),     //            .writedata
		.avalon_readdata      (mm_interconnect_0_buffered_spi_0_avalon_readdata),      //            .readdata
		.avalon_readdatavalid (mm_interconnect_0_buffered_spi_0_avalon_readdatavalid), //            .readdatavalid
		.spi_mosi             (buffered_spi_mosi),                                     // conduit_end.mosi
		.spi_clk              (buffered_spi_clk),                                      //            .clk
		.spi_miso             (buffered_spi_miso),                                     //            .miso
		.spi_cs               (buffered_spi_cs),                                       //            .cs
		.clock                (clock_116_mhz_clk)                                      //       clock.clk
	);

	wasca_extra_leds extra_leds (
		.clk        (clock_116_mhz_clk),                          //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_extra_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_extra_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_extra_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_extra_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_extra_leds_s1_readdata),   //                    .readdata
		.out_port   (extra_leds_conn_export)                      // external_connection.export
	);

	wasca_hex0 hex0 (
		.clk        (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_hex0_s1_address),       //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_s1_write),        //                    .write_n
		.writedata  (mm_interconnect_0_hex0_s1_writedata),     //                    .writedata
		.chipselect (mm_interconnect_0_hex0_s1_chipselect),    //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_s1_readdata),      //                    .readdata
		.out_port   (hex0_conn_export)                         // external_connection.export
	);

	wasca_hex0 hex1 (
		.clk        (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_hex1_s1_address),       //                  s1.address
		.write_n    (~mm_interconnect_0_hex1_s1_write),        //                    .write_n
		.writedata  (mm_interconnect_0_hex1_s1_writedata),     //                    .writedata
		.chipselect (mm_interconnect_0_hex1_s1_chipselect),    //                    .chipselect
		.readdata   (mm_interconnect_0_hex1_s1_readdata),      //                    .readdata
		.out_port   (hex1_conn_export)                         // external_connection.export
	);

	wasca_hex0 hex2 (
		.clk        (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_hex2_s1_address),       //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_s1_write),        //                    .write_n
		.writedata  (mm_interconnect_0_hex2_s1_writedata),     //                    .writedata
		.chipselect (mm_interconnect_0_hex2_s1_chipselect),    //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_s1_readdata),      //                    .readdata
		.out_port   (hex2_conn_export)                         // external_connection.export
	);

	wasca_hex0 hex3 (
		.clk        (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_hex3_s1_address),       //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_s1_write),        //                    .write_n
		.writedata  (mm_interconnect_0_hex3_s1_writedata),     //                    .writedata
		.chipselect (mm_interconnect_0_hex3_s1_chipselect),    //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_s1_readdata),      //                    .readdata
		.out_port   (hex3_conn_export)                         // external_connection.export
	);

	wasca_hex0 hex4 (
		.clk        (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_hex4_s1_address),       //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_s1_write),        //                    .write_n
		.writedata  (mm_interconnect_0_hex4_s1_writedata),     //                    .writedata
		.chipselect (mm_interconnect_0_hex4_s1_chipselect),    //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_s1_readdata),      //                    .readdata
		.out_port   (hex4_conn_export)                         // external_connection.export
	);

	wasca_hex0 hex5 (
		.clk        (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_hex5_s1_address),       //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_s1_write),        //                    .write_n
		.writedata  (mm_interconnect_0_hex5_s1_writedata),     //                    .writedata
		.chipselect (mm_interconnect_0_hex5_s1_chipselect),    //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_s1_readdata),      //                    .readdata
		.out_port   (hex5_conn_export)                         // external_connection.export
	);

	wasca_hexdot hexdot (
		.clk        (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_hexdot_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_0_hexdot_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_0_hexdot_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_0_hexdot_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_0_hexdot_s1_readdata),    //                    .readdata
		.out_port   (hexdot_conn_export)                       // external_connection.export
	);

	wasca_leds leds (
		.clk        (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n    (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),       //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),        //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),     //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect),    //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),      //                    .readdata
		.out_port   (leds_conn_export)                         // external_connection.export
	);

	wasca_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clock_116_mhz_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M50DAF484C7G"),
		.DEVICE_ID                           ("50"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (8191),
		.SECTOR2_START_ADDR                  (8192),
		.SECTOR2_END_ADDR                    (16383),
		.SECTOR3_START_ADDR                  (16384),
		.SECTOR3_END_ADDR                    (114687),
		.SECTOR4_START_ADDR                  (114688),
		.SECTOR4_END_ADDR                    (188415),
		.SECTOR5_START_ADDR                  (188416),
		.SECTOR5_END_ADDR                    (360447),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (360447),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (114687),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (360447),
		.ADDR_RANGE1_OFFSET                  (2048),
		.ADDR_RANGE2_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (19),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (0),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (5),
		.FLASH_RESET_CYCLE_MAX_INDEX         (29),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (139),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (40603248),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (35382),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("False")
	) onchip_flash_0 (
		.clock                   (clock_116_mhz_clk),                                   //    clk.clk
		.reset_n                 (~rst_controller_reset_out_reset),                     // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_onchip_flash_0_csr_readdata)        //       .readdata
	);

	wasca_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clock_116_mhz_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	wasca_performance_counter_0 performance_counter_0 (
		.clk           (clock_116_mhz_clk),                                                   //           clk.clk
		.reset_n       (~nios2_gen2_0_debug_reset_request_reset),                             //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_0_control_slave_writedata)      //              .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_0 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (reset_controller_0_reset_in1_reset),     // reset_in1.reset
		.clk            (clock_116_mhz_clk),                      //       clk.clk
		.reset_out      (reset_controller_0_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	wasca_spi_sync spi_sync (
		.clk      (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n  (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address  (mm_interconnect_0_spi_sync_s1_address),   //                  s1.address
		.readdata (mm_interconnect_0_spi_sync_s1_readdata),  //                    .readdata
		.in_port  (spi_sync_conn_export)                     // external_connection.export
	);

	wasca_switches switches (
		.clk      (clock_116_mhz_clk),                       //                 clk.clk
		.reset_n  (~nios2_gen2_0_debug_reset_request_reset), //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),   //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata),  //                    .readdata
		.in_port  (switches_conn_export)                     // external_connection.export
	);

	wasca_uart_0 uart_0 (
		.clk           (clock_116_mhz_clk),                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.dataavailable (),                                          //                    .dataavailable
		.readyfordata  (),                                          //                    .readyfordata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver0_irq)                   //                 irq.irq
	);

	wasca_mm_interconnect_0 mm_interconnect_0 (
		.altpll_1_c0_clk                                            (clock_116_mhz_clk),                                                       //                                          altpll_1_c0.clk
		.clk_0_clk_clk                                              (clk_clk),                                                                 //                                            clk_0_clk.clk
		.altpll_1_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                      // altpll_1_inclk_interface_reset_reset_bridge_in_reset.reset
		.buffered_spi_0_reset_reset_bridge_in_reset_reset           (nios2_gen2_0_debug_reset_request_reset),                                  //           buffered_spi_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                          //             nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                           (nios2_gen2_0_data_master_address),                                        //                             nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                                    //                                                     .waitrequest
		.nios2_gen2_0_data_master_byteenable                        (nios2_gen2_0_data_master_byteenable),                                     //                                                     .byteenable
		.nios2_gen2_0_data_master_read                              (nios2_gen2_0_data_master_read),                                           //                                                     .read
		.nios2_gen2_0_data_master_readdata                          (nios2_gen2_0_data_master_readdata),                                       //                                                     .readdata
		.nios2_gen2_0_data_master_write                             (nios2_gen2_0_data_master_write),                                          //                                                     .write
		.nios2_gen2_0_data_master_writedata                         (nios2_gen2_0_data_master_writedata),                                      //                                                     .writedata
		.nios2_gen2_0_data_master_debugaccess                       (nios2_gen2_0_data_master_debugaccess),                                    //                                                     .debugaccess
		.nios2_gen2_0_instruction_master_address                    (nios2_gen2_0_instruction_master_address),                                 //                      nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                (nios2_gen2_0_instruction_master_waitrequest),                             //                                                     .waitrequest
		.nios2_gen2_0_instruction_master_read                       (nios2_gen2_0_instruction_master_read),                                    //                                                     .read
		.nios2_gen2_0_instruction_master_readdata                   (nios2_gen2_0_instruction_master_readdata),                                //                                                     .readdata
		.abus_avalon_sdram_bridge_0_avalon_regs_address             (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_address),        //               abus_avalon_sdram_bridge_0_avalon_regs.address
		.abus_avalon_sdram_bridge_0_avalon_regs_write               (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_write),          //                                                     .write
		.abus_avalon_sdram_bridge_0_avalon_regs_read                (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_read),           //                                                     .read
		.abus_avalon_sdram_bridge_0_avalon_regs_readdata            (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_readdata),       //                                                     .readdata
		.abus_avalon_sdram_bridge_0_avalon_regs_writedata           (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_writedata),      //                                                     .writedata
		.abus_avalon_sdram_bridge_0_avalon_regs_readdatavalid       (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_readdatavalid),  //                                                     .readdatavalid
		.abus_avalon_sdram_bridge_0_avalon_regs_waitrequest         (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_regs_waitrequest),    //                                                     .waitrequest
		.abus_avalon_sdram_bridge_0_avalon_sdram_address            (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_address),       //              abus_avalon_sdram_bridge_0_avalon_sdram.address
		.abus_avalon_sdram_bridge_0_avalon_sdram_write              (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_write),         //                                                     .write
		.abus_avalon_sdram_bridge_0_avalon_sdram_read               (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_read),          //                                                     .read
		.abus_avalon_sdram_bridge_0_avalon_sdram_readdata           (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_readdata),      //                                                     .readdata
		.abus_avalon_sdram_bridge_0_avalon_sdram_writedata          (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_writedata),     //                                                     .writedata
		.abus_avalon_sdram_bridge_0_avalon_sdram_byteenable         (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_byteenable),    //                                                     .byteenable
		.abus_avalon_sdram_bridge_0_avalon_sdram_readdatavalid      (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_readdatavalid), //                                                     .readdatavalid
		.abus_avalon_sdram_bridge_0_avalon_sdram_waitrequest        (mm_interconnect_0_abus_avalon_sdram_bridge_0_avalon_sdram_waitrequest),   //                                                     .waitrequest
		.altpll_1_pll_slave_address                                 (mm_interconnect_0_altpll_1_pll_slave_address),                            //                                   altpll_1_pll_slave.address
		.altpll_1_pll_slave_write                                   (mm_interconnect_0_altpll_1_pll_slave_write),                              //                                                     .write
		.altpll_1_pll_slave_read                                    (mm_interconnect_0_altpll_1_pll_slave_read),                               //                                                     .read
		.altpll_1_pll_slave_readdata                                (mm_interconnect_0_altpll_1_pll_slave_readdata),                           //                                                     .readdata
		.altpll_1_pll_slave_writedata                               (mm_interconnect_0_altpll_1_pll_slave_writedata),                          //                                                     .writedata
		.buffered_spi_0_avalon_address                              (mm_interconnect_0_buffered_spi_0_avalon_address),                         //                                buffered_spi_0_avalon.address
		.buffered_spi_0_avalon_write                                (mm_interconnect_0_buffered_spi_0_avalon_write),                           //                                                     .write
		.buffered_spi_0_avalon_read                                 (mm_interconnect_0_buffered_spi_0_avalon_read),                            //                                                     .read
		.buffered_spi_0_avalon_readdata                             (mm_interconnect_0_buffered_spi_0_avalon_readdata),                        //                                                     .readdata
		.buffered_spi_0_avalon_writedata                            (mm_interconnect_0_buffered_spi_0_avalon_writedata),                       //                                                     .writedata
		.buffered_spi_0_avalon_readdatavalid                        (mm_interconnect_0_buffered_spi_0_avalon_readdatavalid),                   //                                                     .readdatavalid
		.buffered_spi_0_avalon_waitrequest                          (mm_interconnect_0_buffered_spi_0_avalon_waitrequest),                     //                                                     .waitrequest
		.extra_leds_s1_address                                      (mm_interconnect_0_extra_leds_s1_address),                                 //                                        extra_leds_s1.address
		.extra_leds_s1_write                                        (mm_interconnect_0_extra_leds_s1_write),                                   //                                                     .write
		.extra_leds_s1_readdata                                     (mm_interconnect_0_extra_leds_s1_readdata),                                //                                                     .readdata
		.extra_leds_s1_writedata                                    (mm_interconnect_0_extra_leds_s1_writedata),                               //                                                     .writedata
		.extra_leds_s1_chipselect                                   (mm_interconnect_0_extra_leds_s1_chipselect),                              //                                                     .chipselect
		.hex0_s1_address                                            (mm_interconnect_0_hex0_s1_address),                                       //                                              hex0_s1.address
		.hex0_s1_write                                              (mm_interconnect_0_hex0_s1_write),                                         //                                                     .write
		.hex0_s1_readdata                                           (mm_interconnect_0_hex0_s1_readdata),                                      //                                                     .readdata
		.hex0_s1_writedata                                          (mm_interconnect_0_hex0_s1_writedata),                                     //                                                     .writedata
		.hex0_s1_chipselect                                         (mm_interconnect_0_hex0_s1_chipselect),                                    //                                                     .chipselect
		.hex1_s1_address                                            (mm_interconnect_0_hex1_s1_address),                                       //                                              hex1_s1.address
		.hex1_s1_write                                              (mm_interconnect_0_hex1_s1_write),                                         //                                                     .write
		.hex1_s1_readdata                                           (mm_interconnect_0_hex1_s1_readdata),                                      //                                                     .readdata
		.hex1_s1_writedata                                          (mm_interconnect_0_hex1_s1_writedata),                                     //                                                     .writedata
		.hex1_s1_chipselect                                         (mm_interconnect_0_hex1_s1_chipselect),                                    //                                                     .chipselect
		.hex2_s1_address                                            (mm_interconnect_0_hex2_s1_address),                                       //                                              hex2_s1.address
		.hex2_s1_write                                              (mm_interconnect_0_hex2_s1_write),                                         //                                                     .write
		.hex2_s1_readdata                                           (mm_interconnect_0_hex2_s1_readdata),                                      //                                                     .readdata
		.hex2_s1_writedata                                          (mm_interconnect_0_hex2_s1_writedata),                                     //                                                     .writedata
		.hex2_s1_chipselect                                         (mm_interconnect_0_hex2_s1_chipselect),                                    //                                                     .chipselect
		.hex3_s1_address                                            (mm_interconnect_0_hex3_s1_address),                                       //                                              hex3_s1.address
		.hex3_s1_write                                              (mm_interconnect_0_hex3_s1_write),                                         //                                                     .write
		.hex3_s1_readdata                                           (mm_interconnect_0_hex3_s1_readdata),                                      //                                                     .readdata
		.hex3_s1_writedata                                          (mm_interconnect_0_hex3_s1_writedata),                                     //                                                     .writedata
		.hex3_s1_chipselect                                         (mm_interconnect_0_hex3_s1_chipselect),                                    //                                                     .chipselect
		.hex4_s1_address                                            (mm_interconnect_0_hex4_s1_address),                                       //                                              hex4_s1.address
		.hex4_s1_write                                              (mm_interconnect_0_hex4_s1_write),                                         //                                                     .write
		.hex4_s1_readdata                                           (mm_interconnect_0_hex4_s1_readdata),                                      //                                                     .readdata
		.hex4_s1_writedata                                          (mm_interconnect_0_hex4_s1_writedata),                                     //                                                     .writedata
		.hex4_s1_chipselect                                         (mm_interconnect_0_hex4_s1_chipselect),                                    //                                                     .chipselect
		.hex5_s1_address                                            (mm_interconnect_0_hex5_s1_address),                                       //                                              hex5_s1.address
		.hex5_s1_write                                              (mm_interconnect_0_hex5_s1_write),                                         //                                                     .write
		.hex5_s1_readdata                                           (mm_interconnect_0_hex5_s1_readdata),                                      //                                                     .readdata
		.hex5_s1_writedata                                          (mm_interconnect_0_hex5_s1_writedata),                                     //                                                     .writedata
		.hex5_s1_chipselect                                         (mm_interconnect_0_hex5_s1_chipselect),                                    //                                                     .chipselect
		.hexdot_s1_address                                          (mm_interconnect_0_hexdot_s1_address),                                     //                                            hexdot_s1.address
		.hexdot_s1_write                                            (mm_interconnect_0_hexdot_s1_write),                                       //                                                     .write
		.hexdot_s1_readdata                                         (mm_interconnect_0_hexdot_s1_readdata),                                    //                                                     .readdata
		.hexdot_s1_writedata                                        (mm_interconnect_0_hexdot_s1_writedata),                                   //                                                     .writedata
		.hexdot_s1_chipselect                                       (mm_interconnect_0_hexdot_s1_chipselect),                                  //                                                     .chipselect
		.leds_s1_address                                            (mm_interconnect_0_leds_s1_address),                                       //                                              leds_s1.address
		.leds_s1_write                                              (mm_interconnect_0_leds_s1_write),                                         //                                                     .write
		.leds_s1_readdata                                           (mm_interconnect_0_leds_s1_readdata),                                      //                                                     .readdata
		.leds_s1_writedata                                          (mm_interconnect_0_leds_s1_writedata),                                     //                                                     .writedata
		.leds_s1_chipselect                                         (mm_interconnect_0_leds_s1_chipselect),                                    //                                                     .chipselect
		.nios2_gen2_0_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                  //                         nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                    //                                                     .write
		.nios2_gen2_0_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                     //                                                     .read
		.nios2_gen2_0_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),                 //                                                     .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),                //                                                     .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),               //                                                     .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),              //                                                     .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),              //                                                     .debugaccess
		.onchip_flash_0_csr_address                                 (mm_interconnect_0_onchip_flash_0_csr_address),                            //                                   onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                                   (mm_interconnect_0_onchip_flash_0_csr_write),                              //                                                     .write
		.onchip_flash_0_csr_read                                    (mm_interconnect_0_onchip_flash_0_csr_read),                               //                                                     .read
		.onchip_flash_0_csr_readdata                                (mm_interconnect_0_onchip_flash_0_csr_readdata),                           //                                                     .readdata
		.onchip_flash_0_csr_writedata                               (mm_interconnect_0_onchip_flash_0_csr_writedata),                          //                                                     .writedata
		.onchip_flash_0_data_address                                (mm_interconnect_0_onchip_flash_0_data_address),                           //                                  onchip_flash_0_data.address
		.onchip_flash_0_data_write                                  (mm_interconnect_0_onchip_flash_0_data_write),                             //                                                     .write
		.onchip_flash_0_data_read                                   (mm_interconnect_0_onchip_flash_0_data_read),                              //                                                     .read
		.onchip_flash_0_data_readdata                               (mm_interconnect_0_onchip_flash_0_data_readdata),                          //                                                     .readdata
		.onchip_flash_0_data_writedata                              (mm_interconnect_0_onchip_flash_0_data_writedata),                         //                                                     .writedata
		.onchip_flash_0_data_burstcount                             (mm_interconnect_0_onchip_flash_0_data_burstcount),                        //                                                     .burstcount
		.onchip_flash_0_data_readdatavalid                          (mm_interconnect_0_onchip_flash_0_data_readdatavalid),                     //                                                     .readdatavalid
		.onchip_flash_0_data_waitrequest                            (mm_interconnect_0_onchip_flash_0_data_waitrequest),                       //                                                     .waitrequest
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                           //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                             //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),                          //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),                         //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                        //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                        //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                             //                                                     .clken
		.performance_counter_0_control_slave_address                (mm_interconnect_0_performance_counter_0_control_slave_address),           //                  performance_counter_0_control_slave.address
		.performance_counter_0_control_slave_write                  (mm_interconnect_0_performance_counter_0_control_slave_write),             //                                                     .write
		.performance_counter_0_control_slave_readdata               (mm_interconnect_0_performance_counter_0_control_slave_readdata),          //                                                     .readdata
		.performance_counter_0_control_slave_writedata              (mm_interconnect_0_performance_counter_0_control_slave_writedata),         //                                                     .writedata
		.performance_counter_0_control_slave_begintransfer          (mm_interconnect_0_performance_counter_0_control_slave_begintransfer),     //                                                     .begintransfer
		.spi_sync_s1_address                                        (mm_interconnect_0_spi_sync_s1_address),                                   //                                          spi_sync_s1.address
		.spi_sync_s1_readdata                                       (mm_interconnect_0_spi_sync_s1_readdata),                                  //                                                     .readdata
		.switches_s1_address                                        (mm_interconnect_0_switches_s1_address),                                   //                                          switches_s1.address
		.switches_s1_readdata                                       (mm_interconnect_0_switches_s1_readdata),                                  //                                                     .readdata
		.uart_0_s1_address                                          (mm_interconnect_0_uart_0_s1_address),                                     //                                            uart_0_s1.address
		.uart_0_s1_write                                            (mm_interconnect_0_uart_0_s1_write),                                       //                                                     .write
		.uart_0_s1_read                                             (mm_interconnect_0_uart_0_s1_read),                                        //                                                     .read
		.uart_0_s1_readdata                                         (mm_interconnect_0_uart_0_s1_readdata),                                    //                                                     .readdata
		.uart_0_s1_writedata                                        (mm_interconnect_0_uart_0_s1_writedata),                                   //                                                     .writedata
		.uart_0_s1_begintransfer                                    (mm_interconnect_0_uart_0_s1_begintransfer),                               //                                                     .begintransfer
		.uart_0_s1_chipselect                                       (mm_interconnect_0_uart_0_s1_chipselect)                                   //                                                     .chipselect
	);

	wasca_irq_mapper irq_mapper (
		.clk           (clock_116_mhz_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_controller_0_reset_out_reset), // reset_in0.reset
		.clk            (clock_116_mhz_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (reset_controller_0_reset_out_reset), // reset_in0.reset
		.clk            (clock_116_mhz_clk),                  //       clk.clk
		.reset_out      (),                                   // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
