// wasca.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module wasca (
		input  wire [9:0]  abus_slave_0_abus_address,                      //                 abus_slave_0_abus.address
		input  wire [2:0]  abus_slave_0_abus_chipselect,                   //                                  .chipselect
		input  wire        abus_slave_0_abus_read,                         //                                  .read
		input  wire [1:0]  abus_slave_0_abus_write,                        //                                  .write
		output wire        abus_slave_0_abus_waitrequest,                  //                                  .waitrequest
		output wire        abus_slave_0_abus_interrupt,                    //                                  .interrupt
		inout  wire [15:0] abus_slave_0_abus_addressdata,                  //                                  .addressdata
		output wire        abus_slave_0_abus_direction,                    //                                  .direction
		output wire [1:0]  abus_slave_0_abus_muxing,                       //                                  .muxing
		output wire        abus_slave_0_abus_disableout,                   //                                  .disableout
		input  wire        abus_slave_0_conduit_saturn_reset_saturn_reset, // abus_slave_0_conduit_saturn_reset.saturn_reset
		input  wire        altpll_0_areset_conduit_export,                 //           altpll_0_areset_conduit.export
		output wire        altpll_0_locked_conduit_export,                 //           altpll_0_locked_conduit.export
		output wire        altpll_0_phasedone_conduit_export,              //        altpll_0_phasedone_conduit.export
		input  wire        clk_clk,                                        //                               clk.clk
		output wire [12:0] external_sdram_controller_wire_addr,            //    external_sdram_controller_wire.addr
		output wire [1:0]  external_sdram_controller_wire_ba,              //                                  .ba
		output wire        external_sdram_controller_wire_cas_n,           //                                  .cas_n
		output wire        external_sdram_controller_wire_cke,             //                                  .cke
		output wire        external_sdram_controller_wire_cs_n,            //                                  .cs_n
		inout  wire [15:0] external_sdram_controller_wire_dq,              //                                  .dq
		output wire [1:0]  external_sdram_controller_wire_dqm,             //                                  .dqm
		output wire        external_sdram_controller_wire_ras_n,           //                                  .ras_n
		output wire        external_sdram_controller_wire_we_n,            //                                  .we_n
		output wire [4:0]  extra_leds_conn_export,                         //                   extra_leds_conn.export
		output wire [6:0]  hex0_conn_export,                               //                         hex0_conn.export
		output wire [6:0]  hex1_conn_export,                               //                         hex1_conn.export
		output wire [6:0]  hex2_conn_export,                               //                         hex2_conn.export
		output wire [6:0]  hex3_conn_export,                               //                         hex3_conn.export
		output wire [6:0]  hex4_conn_export,                               //                         hex4_conn.export
		output wire [6:0]  hex5_conn_export,                               //                         hex5_conn.export
		output wire [5:0]  hexdot_conn_export,                             //                       hexdot_conn.export
		output wire [3:0]  leds_conn_export,                               //                         leds_conn.export
		output wire        sdram_clkout_clk,                               //                      sdram_clkout.clk
		input  wire        spi_stm32_MISO,                                 //                         spi_stm32.MISO
		output wire        spi_stm32_MOSI,                                 //                                  .MOSI
		output wire        spi_stm32_SCLK,                                 //                                  .SCLK
		output wire        spi_stm32_SS_n,                                 //                                  .SS_n
		input  wire        spi_sync_conn_export,                           //                     spi_sync_conn.export
		input  wire [7:0]  switches_conn_export,                           //                     switches_conn.export
		input  wire        uart_0_external_connection_rxd,                 //        uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd                  //                                  .txd
	);

	wire         altpll_0_c0_clk;                                                     // altpll_0:c0 -> [abus_demux_0:clock, abus_slave_0:clock, external_sdram_controller:clk, extra_leds:clk, hex0:clk, hex1:clk, hex2:clk, hex3:clk, hex4:clk, hex5:clk, hexdot:clk, irq_mapper:clk, leds:clk, mm_interconnect_0:altpll_0_c0_clk, mm_interconnect_1:altpll_0_c0_clk, nios2_gen2_0:clk, onchip_flash_0:clock, onchip_memory2_0:clk, onchip_memory2_1:clk, onchip_trace_mem:clk, performance_counter_0:clk, rst_controller:clk, spi_stm32:clk, spi_sync:clk, switches:clk, uart_0:clk]
	wire  [15:0] abus_slave_0_demux_readdata;                                         // abus_slave_0:demux_readdata -> abus_demux_0:demux_readdata
	wire         abus_demux_0_demux_readpulse;                                        // abus_demux_0:demux_readpulse -> abus_slave_0:demux_readpulse
	wire  [27:0] abus_demux_0_demux_readaddress;                                      // abus_demux_0:demux_readaddress -> abus_slave_0:demux_readaddress
	wire  [15:0] abus_demux_0_demux_data;                                             // abus_demux_0:demux_writedata -> abus_slave_0:demux_writedata
	wire         abus_slave_0_demux_readdatavalid;                                    // abus_slave_0:demux_readdatavalid -> abus_demux_0:demux_readdatavalid
	wire   [1:0] abus_demux_0_demux_write_byteenable;                                 // abus_demux_0:demux_write_byteenable -> abus_slave_0:demux_write_byteenable
	wire  [27:0] abus_demux_0_demux_writeaddress;                                     // abus_demux_0:demux_writeaddress -> abus_slave_0:demux_writeaddress
	wire         abus_demux_0_demux_writepulse;                                       // abus_demux_0:demux_writepulse -> abus_slave_0:demux_writepulse
	wire         nios2_gen2_0_debug_reset_request_reset;                              // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire         abus_slave_0_avalon_master_waitrequest;                              // mm_interconnect_0:abus_slave_0_avalon_master_waitrequest -> abus_slave_0:avalon_waitrequest
	wire  [15:0] abus_slave_0_avalon_master_readdata;                                 // mm_interconnect_0:abus_slave_0_avalon_master_readdata -> abus_slave_0:avalon_readdata
	wire         abus_slave_0_avalon_master_read;                                     // abus_slave_0:avalon_read -> mm_interconnect_0:abus_slave_0_avalon_master_read
	wire  [27:0] abus_slave_0_avalon_master_address;                                  // abus_slave_0:avalon_address -> mm_interconnect_0:abus_slave_0_avalon_master_address
	wire   [1:0] abus_slave_0_avalon_master_byteenable;                               // abus_slave_0:avalon_byteenable -> mm_interconnect_0:abus_slave_0_avalon_master_byteenable
	wire         abus_slave_0_avalon_master_readdatavalid;                            // mm_interconnect_0:abus_slave_0_avalon_master_readdatavalid -> abus_slave_0:avalon_readdatavalid
	wire         abus_slave_0_avalon_master_write;                                    // abus_slave_0:avalon_write -> mm_interconnect_0:abus_slave_0_avalon_master_write
	wire  [15:0] abus_slave_0_avalon_master_writedata;                                // abus_slave_0:avalon_writedata -> mm_interconnect_0:abus_slave_0_avalon_master_writedata
	wire         abus_slave_0_avalon_master_burstcount;                               // abus_slave_0:avalon_burstcount -> mm_interconnect_0:abus_slave_0_avalon_master_burstcount
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                   // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                                    // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                 // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                       // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                      // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                  // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                            // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                             // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_external_sdram_controller_s1_chipselect;           // mm_interconnect_0:external_sdram_controller_s1_chipselect -> external_sdram_controller:az_cs
	wire  [15:0] mm_interconnect_0_external_sdram_controller_s1_readdata;             // external_sdram_controller:za_data -> mm_interconnect_0:external_sdram_controller_s1_readdata
	wire         mm_interconnect_0_external_sdram_controller_s1_waitrequest;          // external_sdram_controller:za_waitrequest -> mm_interconnect_0:external_sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_external_sdram_controller_s1_address;              // mm_interconnect_0:external_sdram_controller_s1_address -> external_sdram_controller:az_addr
	wire         mm_interconnect_0_external_sdram_controller_s1_read;                 // mm_interconnect_0:external_sdram_controller_s1_read -> external_sdram_controller:az_rd_n
	wire   [1:0] mm_interconnect_0_external_sdram_controller_s1_byteenable;           // mm_interconnect_0:external_sdram_controller_s1_byteenable -> external_sdram_controller:az_be_n
	wire         mm_interconnect_0_external_sdram_controller_s1_readdatavalid;        // external_sdram_controller:za_valid -> mm_interconnect_0:external_sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_external_sdram_controller_s1_write;                // mm_interconnect_0:external_sdram_controller_s1_write -> external_sdram_controller:az_wr_n
	wire  [15:0] mm_interconnect_0_external_sdram_controller_s1_writedata;            // mm_interconnect_0:external_sdram_controller_s1_writedata -> external_sdram_controller:az_data
	wire         mm_interconnect_0_onchip_memory2_1_s1_chipselect;                    // mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_readdata;                      // onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_1_s1_address;                       // mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_1_s1_byteenable;                    // mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	wire         mm_interconnect_0_onchip_memory2_1_s1_write;                         // mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_writedata;                     // mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_clken;                         // mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	wire  [31:0] mm_interconnect_0_abus_slave_0_avalon_nios_readdata;                 // abus_slave_0:avalon_nios_readdata -> mm_interconnect_0:abus_slave_0_avalon_nios_readdata
	wire         mm_interconnect_0_abus_slave_0_avalon_nios_waitrequest;              // abus_slave_0:avalon_nios_waitrequest -> mm_interconnect_0:abus_slave_0_avalon_nios_waitrequest
	wire   [7:0] mm_interconnect_0_abus_slave_0_avalon_nios_address;                  // mm_interconnect_0:abus_slave_0_avalon_nios_address -> abus_slave_0:avalon_nios_address
	wire         mm_interconnect_0_abus_slave_0_avalon_nios_read;                     // mm_interconnect_0:abus_slave_0_avalon_nios_read -> abus_slave_0:avalon_nios_read
	wire         mm_interconnect_0_abus_slave_0_avalon_nios_readdatavalid;            // abus_slave_0:avalon_nios_readdatavalid -> mm_interconnect_0:abus_slave_0_avalon_nios_readdatavalid
	wire         mm_interconnect_0_abus_slave_0_avalon_nios_write;                    // mm_interconnect_0:abus_slave_0_avalon_nios_write -> abus_slave_0:avalon_nios_write
	wire  [31:0] mm_interconnect_0_abus_slave_0_avalon_nios_writedata;                // mm_interconnect_0:abus_slave_0_avalon_nios_writedata -> abus_slave_0:avalon_nios_writedata
	wire   [0:0] mm_interconnect_0_abus_slave_0_avalon_nios_burstcount;               // mm_interconnect_0:abus_slave_0_avalon_nios_burstcount -> abus_slave_0:avalon_nios_burstcount
	wire  [31:0] mm_interconnect_0_abus_demux_0_avalon_nios_readdata;                 // abus_demux_0:avalon_nios_readdata -> mm_interconnect_0:abus_demux_0_avalon_nios_readdata
	wire         mm_interconnect_0_abus_demux_0_avalon_nios_waitrequest;              // abus_demux_0:avalon_nios_waitrequest -> mm_interconnect_0:abus_demux_0_avalon_nios_waitrequest
	wire   [7:0] mm_interconnect_0_abus_demux_0_avalon_nios_address;                  // mm_interconnect_0:abus_demux_0_avalon_nios_address -> abus_demux_0:avalon_nios_address
	wire         mm_interconnect_0_abus_demux_0_avalon_nios_read;                     // mm_interconnect_0:abus_demux_0_avalon_nios_read -> abus_demux_0:avalon_nios_read
	wire         mm_interconnect_0_abus_demux_0_avalon_nios_readdatavalid;            // abus_demux_0:avalon_nios_readdatavalid -> mm_interconnect_0:abus_demux_0_avalon_nios_readdatavalid
	wire         mm_interconnect_0_abus_demux_0_avalon_nios_write;                    // mm_interconnect_0:abus_demux_0_avalon_nios_write -> abus_demux_0:avalon_nios_write
	wire  [31:0] mm_interconnect_0_abus_demux_0_avalon_nios_writedata;                // mm_interconnect_0:abus_demux_0_avalon_nios_writedata -> abus_demux_0:avalon_nios_writedata
	wire   [0:0] mm_interconnect_0_abus_demux_0_avalon_nios_burstcount;               // mm_interconnect_0:abus_demux_0_avalon_nios_burstcount -> abus_demux_0:avalon_nios_burstcount
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_readdata;      // performance_counter_0:readdata -> mm_interconnect_0:performance_counter_0_control_slave_readdata
	wire   [2:0] mm_interconnect_0_performance_counter_0_control_slave_address;       // mm_interconnect_0:performance_counter_0_control_slave_address -> performance_counter_0:address
	wire         mm_interconnect_0_performance_counter_0_control_slave_begintransfer; // mm_interconnect_0:performance_counter_0_control_slave_begintransfer -> performance_counter_0:begintransfer
	wire         mm_interconnect_0_performance_counter_0_control_slave_write;         // mm_interconnect_0:performance_counter_0_control_slave_write -> performance_counter_0:write
	wire  [31:0] mm_interconnect_0_performance_counter_0_control_slave_writedata;     // mm_interconnect_0:performance_counter_0_control_slave_writedata -> performance_counter_0:writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_readdata;                       // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	wire   [0:0] mm_interconnect_0_onchip_flash_0_csr_address;                        // mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_0_onchip_flash_0_csr_read;                           // mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire         mm_interconnect_0_onchip_flash_0_csr_write;                          // mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_writedata;                      // mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;                      // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;                   // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire  [18:0] mm_interconnect_0_onchip_flash_0_data_address;                       // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_read;                          // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;                 // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_onchip_flash_0_data_write;                         // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;                     // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;                    // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;             // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;          // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                 // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                       // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                        // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                           // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                          // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                      // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                    // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                      // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                       // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                    // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                         // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                     // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                         // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                              // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                               // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                  // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                   // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                     // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                 // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                              // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                                // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                 // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                    // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                           // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                   // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                               // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_hex0_s1_chipselect;                                // mm_interconnect_0:hex0_s1_chipselect -> hex0:chipselect
	wire  [31:0] mm_interconnect_0_hex0_s1_readdata;                                  // hex0:readdata -> mm_interconnect_0:hex0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_s1_address;                                   // mm_interconnect_0:hex0_s1_address -> hex0:address
	wire         mm_interconnect_0_hex0_s1_write;                                     // mm_interconnect_0:hex0_s1_write -> hex0:write_n
	wire  [31:0] mm_interconnect_0_hex0_s1_writedata;                                 // mm_interconnect_0:hex0_s1_writedata -> hex0:writedata
	wire         mm_interconnect_0_hex1_s1_chipselect;                                // mm_interconnect_0:hex1_s1_chipselect -> hex1:chipselect
	wire  [31:0] mm_interconnect_0_hex1_s1_readdata;                                  // hex1:readdata -> mm_interconnect_0:hex1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex1_s1_address;                                   // mm_interconnect_0:hex1_s1_address -> hex1:address
	wire         mm_interconnect_0_hex1_s1_write;                                     // mm_interconnect_0:hex1_s1_write -> hex1:write_n
	wire  [31:0] mm_interconnect_0_hex1_s1_writedata;                                 // mm_interconnect_0:hex1_s1_writedata -> hex1:writedata
	wire         mm_interconnect_0_hex2_s1_chipselect;                                // mm_interconnect_0:hex2_s1_chipselect -> hex2:chipselect
	wire  [31:0] mm_interconnect_0_hex2_s1_readdata;                                  // hex2:readdata -> mm_interconnect_0:hex2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex2_s1_address;                                   // mm_interconnect_0:hex2_s1_address -> hex2:address
	wire         mm_interconnect_0_hex2_s1_write;                                     // mm_interconnect_0:hex2_s1_write -> hex2:write_n
	wire  [31:0] mm_interconnect_0_hex2_s1_writedata;                                 // mm_interconnect_0:hex2_s1_writedata -> hex2:writedata
	wire         mm_interconnect_0_hex3_s1_chipselect;                                // mm_interconnect_0:hex3_s1_chipselect -> hex3:chipselect
	wire  [31:0] mm_interconnect_0_hex3_s1_readdata;                                  // hex3:readdata -> mm_interconnect_0:hex3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_s1_address;                                   // mm_interconnect_0:hex3_s1_address -> hex3:address
	wire         mm_interconnect_0_hex3_s1_write;                                     // mm_interconnect_0:hex3_s1_write -> hex3:write_n
	wire  [31:0] mm_interconnect_0_hex3_s1_writedata;                                 // mm_interconnect_0:hex3_s1_writedata -> hex3:writedata
	wire         mm_interconnect_0_hex4_s1_chipselect;                                // mm_interconnect_0:hex4_s1_chipselect -> hex4:chipselect
	wire  [31:0] mm_interconnect_0_hex4_s1_readdata;                                  // hex4:readdata -> mm_interconnect_0:hex4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_s1_address;                                   // mm_interconnect_0:hex4_s1_address -> hex4:address
	wire         mm_interconnect_0_hex4_s1_write;                                     // mm_interconnect_0:hex4_s1_write -> hex4:write_n
	wire  [31:0] mm_interconnect_0_hex4_s1_writedata;                                 // mm_interconnect_0:hex4_s1_writedata -> hex4:writedata
	wire         mm_interconnect_0_hex5_s1_chipselect;                                // mm_interconnect_0:hex5_s1_chipselect -> hex5:chipselect
	wire  [31:0] mm_interconnect_0_hex5_s1_readdata;                                  // hex5:readdata -> mm_interconnect_0:hex5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_s1_address;                                   // mm_interconnect_0:hex5_s1_address -> hex5:address
	wire         mm_interconnect_0_hex5_s1_write;                                     // mm_interconnect_0:hex5_s1_write -> hex5:write_n
	wire  [31:0] mm_interconnect_0_hex5_s1_writedata;                                 // mm_interconnect_0:hex5_s1_writedata -> hex5:writedata
	wire         mm_interconnect_0_hexdot_s1_chipselect;                              // mm_interconnect_0:hexdot_s1_chipselect -> hexdot:chipselect
	wire  [31:0] mm_interconnect_0_hexdot_s1_readdata;                                // hexdot:readdata -> mm_interconnect_0:hexdot_s1_readdata
	wire   [1:0] mm_interconnect_0_hexdot_s1_address;                                 // mm_interconnect_0:hexdot_s1_address -> hexdot:address
	wire         mm_interconnect_0_hexdot_s1_write;                                   // mm_interconnect_0:hexdot_s1_write -> hexdot:write_n
	wire  [31:0] mm_interconnect_0_hexdot_s1_writedata;                               // mm_interconnect_0:hexdot_s1_writedata -> hexdot:writedata
	wire  [31:0] mm_interconnect_0_spi_sync_s1_readdata;                              // spi_sync:readdata -> mm_interconnect_0:spi_sync_s1_readdata
	wire   [1:0] mm_interconnect_0_spi_sync_s1_address;                               // mm_interconnect_0:spi_sync_s1_address -> spi_sync:address
	wire         mm_interconnect_0_extra_leds_s1_chipselect;                          // mm_interconnect_0:extra_leds_s1_chipselect -> extra_leds:chipselect
	wire  [31:0] mm_interconnect_0_extra_leds_s1_readdata;                            // extra_leds:readdata -> mm_interconnect_0:extra_leds_s1_readdata
	wire   [1:0] mm_interconnect_0_extra_leds_s1_address;                             // mm_interconnect_0:extra_leds_s1_address -> extra_leds:address
	wire         mm_interconnect_0_extra_leds_s1_write;                               // mm_interconnect_0:extra_leds_s1_write -> extra_leds:write_n
	wire  [31:0] mm_interconnect_0_extra_leds_s1_writedata;                           // mm_interconnect_0:extra_leds_s1_writedata -> extra_leds:writedata
	wire         mm_interconnect_0_spi_stm32_spi_control_port_chipselect;             // mm_interconnect_0:spi_stm32_spi_control_port_chipselect -> spi_stm32:spi_select
	wire  [15:0] mm_interconnect_0_spi_stm32_spi_control_port_readdata;               // spi_stm32:data_to_cpu -> mm_interconnect_0:spi_stm32_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_stm32_spi_control_port_address;                // mm_interconnect_0:spi_stm32_spi_control_port_address -> spi_stm32:mem_addr
	wire         mm_interconnect_0_spi_stm32_spi_control_port_read;                   // mm_interconnect_0:spi_stm32_spi_control_port_read -> spi_stm32:read_n
	wire         mm_interconnect_0_spi_stm32_spi_control_port_write;                  // mm_interconnect_0:spi_stm32_spi_control_port_write -> spi_stm32:write_n
	wire  [15:0] mm_interconnect_0_spi_stm32_spi_control_port_writedata;              // mm_interconnect_0:spi_stm32_spi_control_port_writedata -> spi_stm32:data_from_cpu
	wire  [63:0] abus_slave_0_avalon_trace_readdata;                                  // mm_interconnect_1:abus_slave_0_avalon_trace_readdata -> abus_slave_0:avalon_trace_readdata
	wire         abus_slave_0_avalon_trace_waitrequest;                               // mm_interconnect_1:abus_slave_0_avalon_trace_waitrequest -> abus_slave_0:avalon_trace_waitrequest
	wire  [27:0] abus_slave_0_avalon_trace_address;                                   // abus_slave_0:avalon_trace_address -> mm_interconnect_1:abus_slave_0_avalon_trace_address
	wire   [7:0] abus_slave_0_avalon_trace_byteenable;                                // abus_slave_0:avalon_trace_byteenable -> mm_interconnect_1:abus_slave_0_avalon_trace_byteenable
	wire         abus_slave_0_avalon_trace_read;                                      // abus_slave_0:avalon_trace_read -> mm_interconnect_1:abus_slave_0_avalon_trace_read
	wire         abus_slave_0_avalon_trace_readdatavalid;                             // mm_interconnect_1:abus_slave_0_avalon_trace_readdatavalid -> abus_slave_0:avalon_trace_readdatavalid
	wire         abus_slave_0_avalon_trace_write;                                     // abus_slave_0:avalon_trace_write -> mm_interconnect_1:abus_slave_0_avalon_trace_write
	wire  [63:0] abus_slave_0_avalon_trace_writedata;                                 // abus_slave_0:avalon_trace_writedata -> mm_interconnect_1:abus_slave_0_avalon_trace_writedata
	wire         abus_slave_0_avalon_trace_burstcount;                                // abus_slave_0:avalon_trace_burstcount -> mm_interconnect_1:abus_slave_0_avalon_trace_burstcount
	wire         mm_interconnect_1_onchip_trace_mem_s1_chipselect;                    // mm_interconnect_1:onchip_trace_mem_s1_chipselect -> onchip_trace_mem:chipselect
	wire  [63:0] mm_interconnect_1_onchip_trace_mem_s1_readdata;                      // onchip_trace_mem:readdata -> mm_interconnect_1:onchip_trace_mem_s1_readdata
	wire   [8:0] mm_interconnect_1_onchip_trace_mem_s1_address;                       // mm_interconnect_1:onchip_trace_mem_s1_address -> onchip_trace_mem:address
	wire   [7:0] mm_interconnect_1_onchip_trace_mem_s1_byteenable;                    // mm_interconnect_1:onchip_trace_mem_s1_byteenable -> onchip_trace_mem:byteenable
	wire         mm_interconnect_1_onchip_trace_mem_s1_write;                         // mm_interconnect_1:onchip_trace_mem_s1_write -> onchip_trace_mem:write
	wire  [63:0] mm_interconnect_1_onchip_trace_mem_s1_writedata;                     // mm_interconnect_1:onchip_trace_mem_s1_writedata -> onchip_trace_mem:writedata
	wire         mm_interconnect_1_onchip_trace_mem_s1_clken;                         // mm_interconnect_1:onchip_trace_mem_s1_clken -> onchip_trace_mem:clken
	wire         irq_mapper_receiver0_irq;                                            // uart_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                            // spi_stm32:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [abus_demux_0:reset, abus_slave_0:reset, external_sdram_controller:reset_n, extra_leds:reset_n, hex0:reset_n, hex1:reset_n, hex2:reset_n, hex3:reset_n, hex4:reset_n, hex5:reset_n, hexdot:reset_n, irq_mapper:reset, leds:reset_n, mm_interconnect_0:abus_slave_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:abus_slave_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_flash_0:reset_n, onchip_memory2_0:reset, onchip_memory2_1:reset, onchip_trace_mem:reset, performance_counter_0:reset_n, rst_translator:in_reset, spi_stm32:reset_n, spi_sync:reset_n, switches:reset_n, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [onchip_memory2_0:reset_req, onchip_memory2_1:reset_req, onchip_trace_mem:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]

	abus_demux abus_demux_0 (
		.clock                     (altpll_0_c0_clk),                                          //                clock.clk
		.abus_address              (abus_slave_0_abus_address),                                //                 abus.address
		.abus_chipselect           (abus_slave_0_abus_chipselect),                             //                     .chipselect
		.abus_read                 (abus_slave_0_abus_read),                                   //                     .read
		.abus_write                (abus_slave_0_abus_write),                                  //                     .write
		.abus_waitrequest          (abus_slave_0_abus_waitrequest),                            //                     .waitrequest
		.abus_interrupt            (abus_slave_0_abus_interrupt),                              //                     .interrupt
		.abus_addressdata          (abus_slave_0_abus_addressdata),                            //                     .addressdata
		.abus_direction            (abus_slave_0_abus_direction),                              //                     .direction
		.abus_muxing               (abus_slave_0_abus_muxing),                                 //                     .muxing
		.abus_disable_out          (abus_slave_0_abus_disableout),                             //                     .disableout
		.reset                     (rst_controller_reset_out_reset),                           //                reset.reset
		.avalon_nios_read          (mm_interconnect_0_abus_demux_0_avalon_nios_read),          //          avalon_nios.read
		.avalon_nios_write         (mm_interconnect_0_abus_demux_0_avalon_nios_write),         //                     .write
		.avalon_nios_address       (mm_interconnect_0_abus_demux_0_avalon_nios_address),       //                     .address
		.avalon_nios_writedata     (mm_interconnect_0_abus_demux_0_avalon_nios_writedata),     //                     .writedata
		.avalon_nios_readdata      (mm_interconnect_0_abus_demux_0_avalon_nios_readdata),      //                     .readdata
		.avalon_nios_waitrequest   (mm_interconnect_0_abus_demux_0_avalon_nios_waitrequest),   //                     .waitrequest
		.avalon_nios_readdatavalid (mm_interconnect_0_abus_demux_0_avalon_nios_readdatavalid), //                     .readdatavalid
		.avalon_nios_burstcount    (mm_interconnect_0_abus_demux_0_avalon_nios_burstcount),    //                     .burstcount
		.demux_writeaddress        (abus_demux_0_demux_writeaddress),                          //                demux.writeaddress
		.demux_writedata           (abus_demux_0_demux_data),                                  //                     .data
		.demux_writepulse          (abus_demux_0_demux_writepulse),                            //                     .writepulse
		.demux_write_byteenable    (abus_demux_0_demux_write_byteenable),                      //                     .write_byteenable
		.demux_readdata            (abus_slave_0_demux_readdata),                              //                     .readdata
		.demux_readpulse           (abus_demux_0_demux_readpulse),                             //                     .readpulse
		.demux_readdatavalid       (abus_slave_0_demux_readdatavalid),                         //                     .readdatavalid
		.demux_readaddress         (abus_demux_0_demux_readaddress),                           //                     .readaddress
		.saturn_reset              (abus_slave_0_conduit_saturn_reset_saturn_reset)            // conduit_saturn_reset.saturn_reset
	);

	abus_slave abus_slave_0 (
		.clock                      (altpll_0_c0_clk),                                          //         clock.clk
		.avalon_read                (abus_slave_0_avalon_master_read),                          // avalon_master.read
		.avalon_write               (abus_slave_0_avalon_master_write),                         //              .write
		.avalon_waitrequest         (abus_slave_0_avalon_master_waitrequest),                   //              .waitrequest
		.avalon_address             (abus_slave_0_avalon_master_address),                       //              .address
		.avalon_readdata            (abus_slave_0_avalon_master_readdata),                      //              .readdata
		.avalon_writedata           (abus_slave_0_avalon_master_writedata),                     //              .writedata
		.avalon_readdatavalid       (abus_slave_0_avalon_master_readdatavalid),                 //              .readdatavalid
		.avalon_burstcount          (abus_slave_0_avalon_master_burstcount),                    //              .burstcount
		.avalon_byteenable          (abus_slave_0_avalon_master_byteenable),                    //              .byteenable
		.reset                      (rst_controller_reset_out_reset),                           //         reset.reset
		.avalon_nios_read           (mm_interconnect_0_abus_slave_0_avalon_nios_read),          //   avalon_nios.read
		.avalon_nios_write          (mm_interconnect_0_abus_slave_0_avalon_nios_write),         //              .write
		.avalon_nios_address        (mm_interconnect_0_abus_slave_0_avalon_nios_address),       //              .address
		.avalon_nios_writedata      (mm_interconnect_0_abus_slave_0_avalon_nios_writedata),     //              .writedata
		.avalon_nios_readdata       (mm_interconnect_0_abus_slave_0_avalon_nios_readdata),      //              .readdata
		.avalon_nios_waitrequest    (mm_interconnect_0_abus_slave_0_avalon_nios_waitrequest),   //              .waitrequest
		.avalon_nios_readdatavalid  (mm_interconnect_0_abus_slave_0_avalon_nios_readdatavalid), //              .readdatavalid
		.avalon_nios_burstcount     (mm_interconnect_0_abus_slave_0_avalon_nios_burstcount),    //              .burstcount
		.demux_writeaddress         (abus_demux_0_demux_writeaddress),                          //         demux.writeaddress
		.demux_writedata            (abus_demux_0_demux_data),                                  //              .data
		.demux_writepulse           (abus_demux_0_demux_writepulse),                            //              .writepulse
		.demux_write_byteenable     (abus_demux_0_demux_write_byteenable),                      //              .write_byteenable
		.demux_readdata             (abus_slave_0_demux_readdata),                              //              .readdata
		.demux_readpulse            (abus_demux_0_demux_readpulse),                             //              .readpulse
		.demux_readdatavalid        (abus_slave_0_demux_readdatavalid),                         //              .readdatavalid
		.demux_readaddress          (abus_demux_0_demux_readaddress),                           //              .readaddress
		.avalon_trace_address       (abus_slave_0_avalon_trace_address),                        //  avalon_trace.address
		.avalon_trace_burstcount    (abus_slave_0_avalon_trace_burstcount),                     //              .burstcount
		.avalon_trace_byteenable    (abus_slave_0_avalon_trace_byteenable),                     //              .byteenable
		.avalon_trace_read          (abus_slave_0_avalon_trace_read),                           //              .read
		.avalon_trace_readdata      (abus_slave_0_avalon_trace_readdata),                       //              .readdata
		.avalon_trace_readdatavalid (abus_slave_0_avalon_trace_readdatavalid),                  //              .readdatavalid
		.avalon_trace_waitrequest   (abus_slave_0_avalon_trace_waitrequest),                    //              .waitrequest
		.avalon_trace_write         (abus_slave_0_avalon_trace_write),                          //              .write
		.avalon_trace_writedata     (abus_slave_0_avalon_trace_writedata)                       //              .writedata
	);

	wasca_altpll_0 altpll_0 (
		.clk       (clk_clk),                                        //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0        (altpll_0_c0_clk),                                //                    c0.clk
		.c1        (sdram_clkout_clk),                               //                    c1.clk
		.areset    (altpll_0_areset_conduit_export),                 //        areset_conduit.export
		.locked    (altpll_0_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_0_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	wasca_external_sdram_controller external_sdram_controller (
		.clk            (altpll_0_c0_clk),                                              //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                              // reset.reset_n
		.az_addr        (mm_interconnect_0_external_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_external_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_external_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_external_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_external_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_external_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_external_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_external_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_external_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (external_sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (external_sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (external_sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (external_sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (external_sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (external_sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (external_sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (external_sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (external_sdram_controller_wire_we_n)                           //      .export
	);

	wasca_extra_leds extra_leds (
		.clk        (altpll_0_c0_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_extra_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_extra_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_extra_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_extra_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_extra_leds_s1_readdata),   //                    .readdata
		.out_port   (extra_leds_conn_export)                      // external_connection.export
	);

	wasca_hex0 hex0 (
		.clk        (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex0_conn_export)                      // external_connection.export
	);

	wasca_hex0 hex1 (
		.clk        (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex1_s1_readdata),   //                    .readdata
		.out_port   (hex1_conn_export)                      // external_connection.export
	);

	wasca_hex0 hex2 (
		.clk        (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_s1_readdata),   //                    .readdata
		.out_port   (hex2_conn_export)                      // external_connection.export
	);

	wasca_hex0 hex3 (
		.clk        (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_s1_readdata),   //                    .readdata
		.out_port   (hex3_conn_export)                      // external_connection.export
	);

	wasca_hex0 hex4 (
		.clk        (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex4_conn_export)                      // external_connection.export
	);

	wasca_hex0 hex5 (
		.clk        (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_s1_readdata),   //                    .readdata
		.out_port   (hex5_conn_export)                      // external_connection.export
	);

	wasca_hexdot hexdot (
		.clk        (altpll_0_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_hexdot_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hexdot_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hexdot_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hexdot_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hexdot_s1_readdata),   //                    .readdata
		.out_port   (hexdot_conn_export)                      // external_connection.export
	);

	wasca_leds leds (
		.clk        (altpll_0_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_conn_export)                      // external_connection.export
	);

	wasca_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M50DAF484C7G"),
		.DEVICE_ID                           ("50"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (8191),
		.SECTOR2_START_ADDR                  (8192),
		.SECTOR2_END_ADDR                    (16383),
		.SECTOR3_START_ADDR                  (16384),
		.SECTOR3_END_ADDR                    (114687),
		.SECTOR4_START_ADDR                  (114688),
		.SECTOR4_END_ADDR                    (188415),
		.SECTOR5_START_ADDR                  (188416),
		.SECTOR5_END_ADDR                    (360447),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (360447),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (114687),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (360447),
		.ADDR_RANGE1_OFFSET                  (2048),
		.ADDR_RANGE2_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (19),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (0),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (5),
		.FLASH_RESET_CYCLE_MAX_INDEX         (25),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (120),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (35000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (30500),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("False")
	) onchip_flash_0 (
		.clock                   (altpll_0_c0_clk),                                     //    clk.clk
		.reset_n                 (~rst_controller_reset_out_reset),                     // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_onchip_flash_0_csr_readdata)        //       .readdata
	);

	wasca_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	wasca_onchip_memory2_1 onchip_memory2_1 (
		.clk        (altpll_0_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	wasca_onchip_trace_mem onchip_trace_mem (
		.clk        (altpll_0_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_1_onchip_trace_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_trace_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_trace_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_trace_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_trace_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_trace_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_trace_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	wasca_performance_counter_0 performance_counter_0 (
		.clk           (altpll_0_c0_clk),                                                     //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                     //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_0_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_0_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_0_control_slave_writedata)      //              .writedata
	);

	wasca_spi_stm32 spi_stm32 (
		.clk           (altpll_0_c0_clk),                                         //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                         //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_stm32_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_stm32_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_stm32_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_stm32_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_stm32_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_stm32_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver1_irq),                                //              irq.irq
		.MISO          (spi_stm32_MISO),                                          //         external.export
		.MOSI          (spi_stm32_MOSI),                                          //                 .export
		.SCLK          (spi_stm32_SCLK),                                          //                 .export
		.SS_n          (spi_stm32_SS_n)                                           //                 .export
	);

	wasca_spi_sync spi_sync (
		.clk      (altpll_0_c0_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_spi_sync_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_spi_sync_s1_readdata), //                    .readdata
		.in_port  (spi_sync_conn_export)                    // external_connection.export
	);

	wasca_switches switches (
		.clk      (altpll_0_c0_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_conn_export)                    // external_connection.export
	);

	wasca_uart_0 uart_0 (
		.clk           (altpll_0_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.dataavailable (),                                          //                    .dataavailable
		.readyfordata  (),                                          //                    .readyfordata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver0_irq)                   //                 irq.irq
	);

	wasca_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                                     //                                          altpll_0_c0.clk
		.clk_0_clk_clk                                              (clk_clk),                                                             //                                            clk_0_clk.clk
		.abus_slave_0_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                      //             abus_slave_0_reset_reset_bridge_in_reset.reset
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                  // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.abus_slave_0_avalon_master_address                         (abus_slave_0_avalon_master_address),                                  //                           abus_slave_0_avalon_master.address
		.abus_slave_0_avalon_master_waitrequest                     (abus_slave_0_avalon_master_waitrequest),                              //                                                     .waitrequest
		.abus_slave_0_avalon_master_burstcount                      (abus_slave_0_avalon_master_burstcount),                               //                                                     .burstcount
		.abus_slave_0_avalon_master_byteenable                      (abus_slave_0_avalon_master_byteenable),                               //                                                     .byteenable
		.abus_slave_0_avalon_master_read                            (abus_slave_0_avalon_master_read),                                     //                                                     .read
		.abus_slave_0_avalon_master_readdata                        (abus_slave_0_avalon_master_readdata),                                 //                                                     .readdata
		.abus_slave_0_avalon_master_readdatavalid                   (abus_slave_0_avalon_master_readdatavalid),                            //                                                     .readdatavalid
		.abus_slave_0_avalon_master_write                           (abus_slave_0_avalon_master_write),                                    //                                                     .write
		.abus_slave_0_avalon_master_writedata                       (abus_slave_0_avalon_master_writedata),                                //                                                     .writedata
		.nios2_gen2_0_data_master_address                           (nios2_gen2_0_data_master_address),                                    //                             nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                                //                                                     .waitrequest
		.nios2_gen2_0_data_master_byteenable                        (nios2_gen2_0_data_master_byteenable),                                 //                                                     .byteenable
		.nios2_gen2_0_data_master_read                              (nios2_gen2_0_data_master_read),                                       //                                                     .read
		.nios2_gen2_0_data_master_readdata                          (nios2_gen2_0_data_master_readdata),                                   //                                                     .readdata
		.nios2_gen2_0_data_master_write                             (nios2_gen2_0_data_master_write),                                      //                                                     .write
		.nios2_gen2_0_data_master_writedata                         (nios2_gen2_0_data_master_writedata),                                  //                                                     .writedata
		.nios2_gen2_0_data_master_debugaccess                       (nios2_gen2_0_data_master_debugaccess),                                //                                                     .debugaccess
		.nios2_gen2_0_instruction_master_address                    (nios2_gen2_0_instruction_master_address),                             //                      nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                (nios2_gen2_0_instruction_master_waitrequest),                         //                                                     .waitrequest
		.nios2_gen2_0_instruction_master_read                       (nios2_gen2_0_instruction_master_read),                                //                                                     .read
		.nios2_gen2_0_instruction_master_readdata                   (nios2_gen2_0_instruction_master_readdata),                            //                                                     .readdata
		.abus_demux_0_avalon_nios_address                           (mm_interconnect_0_abus_demux_0_avalon_nios_address),                  //                             abus_demux_0_avalon_nios.address
		.abus_demux_0_avalon_nios_write                             (mm_interconnect_0_abus_demux_0_avalon_nios_write),                    //                                                     .write
		.abus_demux_0_avalon_nios_read                              (mm_interconnect_0_abus_demux_0_avalon_nios_read),                     //                                                     .read
		.abus_demux_0_avalon_nios_readdata                          (mm_interconnect_0_abus_demux_0_avalon_nios_readdata),                 //                                                     .readdata
		.abus_demux_0_avalon_nios_writedata                         (mm_interconnect_0_abus_demux_0_avalon_nios_writedata),                //                                                     .writedata
		.abus_demux_0_avalon_nios_burstcount                        (mm_interconnect_0_abus_demux_0_avalon_nios_burstcount),               //                                                     .burstcount
		.abus_demux_0_avalon_nios_readdatavalid                     (mm_interconnect_0_abus_demux_0_avalon_nios_readdatavalid),            //                                                     .readdatavalid
		.abus_demux_0_avalon_nios_waitrequest                       (mm_interconnect_0_abus_demux_0_avalon_nios_waitrequest),              //                                                     .waitrequest
		.abus_slave_0_avalon_nios_address                           (mm_interconnect_0_abus_slave_0_avalon_nios_address),                  //                             abus_slave_0_avalon_nios.address
		.abus_slave_0_avalon_nios_write                             (mm_interconnect_0_abus_slave_0_avalon_nios_write),                    //                                                     .write
		.abus_slave_0_avalon_nios_read                              (mm_interconnect_0_abus_slave_0_avalon_nios_read),                     //                                                     .read
		.abus_slave_0_avalon_nios_readdata                          (mm_interconnect_0_abus_slave_0_avalon_nios_readdata),                 //                                                     .readdata
		.abus_slave_0_avalon_nios_writedata                         (mm_interconnect_0_abus_slave_0_avalon_nios_writedata),                //                                                     .writedata
		.abus_slave_0_avalon_nios_burstcount                        (mm_interconnect_0_abus_slave_0_avalon_nios_burstcount),               //                                                     .burstcount
		.abus_slave_0_avalon_nios_readdatavalid                     (mm_interconnect_0_abus_slave_0_avalon_nios_readdatavalid),            //                                                     .readdatavalid
		.abus_slave_0_avalon_nios_waitrequest                       (mm_interconnect_0_abus_slave_0_avalon_nios_waitrequest),              //                                                     .waitrequest
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                        //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                          //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                           //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                       //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),                      //                                                     .writedata
		.external_sdram_controller_s1_address                       (mm_interconnect_0_external_sdram_controller_s1_address),              //                         external_sdram_controller_s1.address
		.external_sdram_controller_s1_write                         (mm_interconnect_0_external_sdram_controller_s1_write),                //                                                     .write
		.external_sdram_controller_s1_read                          (mm_interconnect_0_external_sdram_controller_s1_read),                 //                                                     .read
		.external_sdram_controller_s1_readdata                      (mm_interconnect_0_external_sdram_controller_s1_readdata),             //                                                     .readdata
		.external_sdram_controller_s1_writedata                     (mm_interconnect_0_external_sdram_controller_s1_writedata),            //                                                     .writedata
		.external_sdram_controller_s1_byteenable                    (mm_interconnect_0_external_sdram_controller_s1_byteenable),           //                                                     .byteenable
		.external_sdram_controller_s1_readdatavalid                 (mm_interconnect_0_external_sdram_controller_s1_readdatavalid),        //                                                     .readdatavalid
		.external_sdram_controller_s1_waitrequest                   (mm_interconnect_0_external_sdram_controller_s1_waitrequest),          //                                                     .waitrequest
		.external_sdram_controller_s1_chipselect                    (mm_interconnect_0_external_sdram_controller_s1_chipselect),           //                                                     .chipselect
		.extra_leds_s1_address                                      (mm_interconnect_0_extra_leds_s1_address),                             //                                        extra_leds_s1.address
		.extra_leds_s1_write                                        (mm_interconnect_0_extra_leds_s1_write),                               //                                                     .write
		.extra_leds_s1_readdata                                     (mm_interconnect_0_extra_leds_s1_readdata),                            //                                                     .readdata
		.extra_leds_s1_writedata                                    (mm_interconnect_0_extra_leds_s1_writedata),                           //                                                     .writedata
		.extra_leds_s1_chipselect                                   (mm_interconnect_0_extra_leds_s1_chipselect),                          //                                                     .chipselect
		.hex0_s1_address                                            (mm_interconnect_0_hex0_s1_address),                                   //                                              hex0_s1.address
		.hex0_s1_write                                              (mm_interconnect_0_hex0_s1_write),                                     //                                                     .write
		.hex0_s1_readdata                                           (mm_interconnect_0_hex0_s1_readdata),                                  //                                                     .readdata
		.hex0_s1_writedata                                          (mm_interconnect_0_hex0_s1_writedata),                                 //                                                     .writedata
		.hex0_s1_chipselect                                         (mm_interconnect_0_hex0_s1_chipselect),                                //                                                     .chipselect
		.hex1_s1_address                                            (mm_interconnect_0_hex1_s1_address),                                   //                                              hex1_s1.address
		.hex1_s1_write                                              (mm_interconnect_0_hex1_s1_write),                                     //                                                     .write
		.hex1_s1_readdata                                           (mm_interconnect_0_hex1_s1_readdata),                                  //                                                     .readdata
		.hex1_s1_writedata                                          (mm_interconnect_0_hex1_s1_writedata),                                 //                                                     .writedata
		.hex1_s1_chipselect                                         (mm_interconnect_0_hex1_s1_chipselect),                                //                                                     .chipselect
		.hex2_s1_address                                            (mm_interconnect_0_hex2_s1_address),                                   //                                              hex2_s1.address
		.hex2_s1_write                                              (mm_interconnect_0_hex2_s1_write),                                     //                                                     .write
		.hex2_s1_readdata                                           (mm_interconnect_0_hex2_s1_readdata),                                  //                                                     .readdata
		.hex2_s1_writedata                                          (mm_interconnect_0_hex2_s1_writedata),                                 //                                                     .writedata
		.hex2_s1_chipselect                                         (mm_interconnect_0_hex2_s1_chipselect),                                //                                                     .chipselect
		.hex3_s1_address                                            (mm_interconnect_0_hex3_s1_address),                                   //                                              hex3_s1.address
		.hex3_s1_write                                              (mm_interconnect_0_hex3_s1_write),                                     //                                                     .write
		.hex3_s1_readdata                                           (mm_interconnect_0_hex3_s1_readdata),                                  //                                                     .readdata
		.hex3_s1_writedata                                          (mm_interconnect_0_hex3_s1_writedata),                                 //                                                     .writedata
		.hex3_s1_chipselect                                         (mm_interconnect_0_hex3_s1_chipselect),                                //                                                     .chipselect
		.hex4_s1_address                                            (mm_interconnect_0_hex4_s1_address),                                   //                                              hex4_s1.address
		.hex4_s1_write                                              (mm_interconnect_0_hex4_s1_write),                                     //                                                     .write
		.hex4_s1_readdata                                           (mm_interconnect_0_hex4_s1_readdata),                                  //                                                     .readdata
		.hex4_s1_writedata                                          (mm_interconnect_0_hex4_s1_writedata),                                 //                                                     .writedata
		.hex4_s1_chipselect                                         (mm_interconnect_0_hex4_s1_chipselect),                                //                                                     .chipselect
		.hex5_s1_address                                            (mm_interconnect_0_hex5_s1_address),                                   //                                              hex5_s1.address
		.hex5_s1_write                                              (mm_interconnect_0_hex5_s1_write),                                     //                                                     .write
		.hex5_s1_readdata                                           (mm_interconnect_0_hex5_s1_readdata),                                  //                                                     .readdata
		.hex5_s1_writedata                                          (mm_interconnect_0_hex5_s1_writedata),                                 //                                                     .writedata
		.hex5_s1_chipselect                                         (mm_interconnect_0_hex5_s1_chipselect),                                //                                                     .chipselect
		.hexdot_s1_address                                          (mm_interconnect_0_hexdot_s1_address),                                 //                                            hexdot_s1.address
		.hexdot_s1_write                                            (mm_interconnect_0_hexdot_s1_write),                                   //                                                     .write
		.hexdot_s1_readdata                                         (mm_interconnect_0_hexdot_s1_readdata),                                //                                                     .readdata
		.hexdot_s1_writedata                                        (mm_interconnect_0_hexdot_s1_writedata),                               //                                                     .writedata
		.hexdot_s1_chipselect                                       (mm_interconnect_0_hexdot_s1_chipselect),                              //                                                     .chipselect
		.leds_s1_address                                            (mm_interconnect_0_leds_s1_address),                                   //                                              leds_s1.address
		.leds_s1_write                                              (mm_interconnect_0_leds_s1_write),                                     //                                                     .write
		.leds_s1_readdata                                           (mm_interconnect_0_leds_s1_readdata),                                  //                                                     .readdata
		.leds_s1_writedata                                          (mm_interconnect_0_leds_s1_writedata),                                 //                                                     .writedata
		.leds_s1_chipselect                                         (mm_interconnect_0_leds_s1_chipselect),                                //                                                     .chipselect
		.nios2_gen2_0_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),              //                         nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                //                                                     .write
		.nios2_gen2_0_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                 //                                                     .read
		.nios2_gen2_0_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),             //                                                     .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),            //                                                     .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),           //                                                     .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),          //                                                     .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),          //                                                     .debugaccess
		.onchip_flash_0_csr_address                                 (mm_interconnect_0_onchip_flash_0_csr_address),                        //                                   onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                                   (mm_interconnect_0_onchip_flash_0_csr_write),                          //                                                     .write
		.onchip_flash_0_csr_read                                    (mm_interconnect_0_onchip_flash_0_csr_read),                           //                                                     .read
		.onchip_flash_0_csr_readdata                                (mm_interconnect_0_onchip_flash_0_csr_readdata),                       //                                                     .readdata
		.onchip_flash_0_csr_writedata                               (mm_interconnect_0_onchip_flash_0_csr_writedata),                      //                                                     .writedata
		.onchip_flash_0_data_address                                (mm_interconnect_0_onchip_flash_0_data_address),                       //                                  onchip_flash_0_data.address
		.onchip_flash_0_data_write                                  (mm_interconnect_0_onchip_flash_0_data_write),                         //                                                     .write
		.onchip_flash_0_data_read                                   (mm_interconnect_0_onchip_flash_0_data_read),                          //                                                     .read
		.onchip_flash_0_data_readdata                               (mm_interconnect_0_onchip_flash_0_data_readdata),                      //                                                     .readdata
		.onchip_flash_0_data_writedata                              (mm_interconnect_0_onchip_flash_0_data_writedata),                     //                                                     .writedata
		.onchip_flash_0_data_burstcount                             (mm_interconnect_0_onchip_flash_0_data_burstcount),                    //                                                     .burstcount
		.onchip_flash_0_data_readdatavalid                          (mm_interconnect_0_onchip_flash_0_data_readdatavalid),                 //                                                     .readdatavalid
		.onchip_flash_0_data_waitrequest                            (mm_interconnect_0_onchip_flash_0_data_waitrequest),                   //                                                     .waitrequest
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                       //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                         //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),                      //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),                     //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                    //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                    //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                         //                                                     .clken
		.onchip_memory2_1_s1_address                                (mm_interconnect_0_onchip_memory2_1_s1_address),                       //                                  onchip_memory2_1_s1.address
		.onchip_memory2_1_s1_write                                  (mm_interconnect_0_onchip_memory2_1_s1_write),                         //                                                     .write
		.onchip_memory2_1_s1_readdata                               (mm_interconnect_0_onchip_memory2_1_s1_readdata),                      //                                                     .readdata
		.onchip_memory2_1_s1_writedata                              (mm_interconnect_0_onchip_memory2_1_s1_writedata),                     //                                                     .writedata
		.onchip_memory2_1_s1_byteenable                             (mm_interconnect_0_onchip_memory2_1_s1_byteenable),                    //                                                     .byteenable
		.onchip_memory2_1_s1_chipselect                             (mm_interconnect_0_onchip_memory2_1_s1_chipselect),                    //                                                     .chipselect
		.onchip_memory2_1_s1_clken                                  (mm_interconnect_0_onchip_memory2_1_s1_clken),                         //                                                     .clken
		.performance_counter_0_control_slave_address                (mm_interconnect_0_performance_counter_0_control_slave_address),       //                  performance_counter_0_control_slave.address
		.performance_counter_0_control_slave_write                  (mm_interconnect_0_performance_counter_0_control_slave_write),         //                                                     .write
		.performance_counter_0_control_slave_readdata               (mm_interconnect_0_performance_counter_0_control_slave_readdata),      //                                                     .readdata
		.performance_counter_0_control_slave_writedata              (mm_interconnect_0_performance_counter_0_control_slave_writedata),     //                                                     .writedata
		.performance_counter_0_control_slave_begintransfer          (mm_interconnect_0_performance_counter_0_control_slave_begintransfer), //                                                     .begintransfer
		.spi_stm32_spi_control_port_address                         (mm_interconnect_0_spi_stm32_spi_control_port_address),                //                           spi_stm32_spi_control_port.address
		.spi_stm32_spi_control_port_write                           (mm_interconnect_0_spi_stm32_spi_control_port_write),                  //                                                     .write
		.spi_stm32_spi_control_port_read                            (mm_interconnect_0_spi_stm32_spi_control_port_read),                   //                                                     .read
		.spi_stm32_spi_control_port_readdata                        (mm_interconnect_0_spi_stm32_spi_control_port_readdata),               //                                                     .readdata
		.spi_stm32_spi_control_port_writedata                       (mm_interconnect_0_spi_stm32_spi_control_port_writedata),              //                                                     .writedata
		.spi_stm32_spi_control_port_chipselect                      (mm_interconnect_0_spi_stm32_spi_control_port_chipselect),             //                                                     .chipselect
		.spi_sync_s1_address                                        (mm_interconnect_0_spi_sync_s1_address),                               //                                          spi_sync_s1.address
		.spi_sync_s1_readdata                                       (mm_interconnect_0_spi_sync_s1_readdata),                              //                                                     .readdata
		.switches_s1_address                                        (mm_interconnect_0_switches_s1_address),                               //                                          switches_s1.address
		.switches_s1_readdata                                       (mm_interconnect_0_switches_s1_readdata),                              //                                                     .readdata
		.uart_0_s1_address                                          (mm_interconnect_0_uart_0_s1_address),                                 //                                            uart_0_s1.address
		.uart_0_s1_write                                            (mm_interconnect_0_uart_0_s1_write),                                   //                                                     .write
		.uart_0_s1_read                                             (mm_interconnect_0_uart_0_s1_read),                                    //                                                     .read
		.uart_0_s1_readdata                                         (mm_interconnect_0_uart_0_s1_readdata),                                //                                                     .readdata
		.uart_0_s1_writedata                                        (mm_interconnect_0_uart_0_s1_writedata),                               //                                                     .writedata
		.uart_0_s1_begintransfer                                    (mm_interconnect_0_uart_0_s1_begintransfer),                           //                                                     .begintransfer
		.uart_0_s1_chipselect                                       (mm_interconnect_0_uart_0_s1_chipselect)                               //                                                     .chipselect
	);

	wasca_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c0_clk                                (altpll_0_c0_clk),                                  //                              altpll_0_c0.clk
		.abus_slave_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // abus_slave_0_reset_reset_bridge_in_reset.reset
		.abus_slave_0_avalon_trace_address              (abus_slave_0_avalon_trace_address),                //                abus_slave_0_avalon_trace.address
		.abus_slave_0_avalon_trace_waitrequest          (abus_slave_0_avalon_trace_waitrequest),            //                                         .waitrequest
		.abus_slave_0_avalon_trace_burstcount           (abus_slave_0_avalon_trace_burstcount),             //                                         .burstcount
		.abus_slave_0_avalon_trace_byteenable           (abus_slave_0_avalon_trace_byteenable),             //                                         .byteenable
		.abus_slave_0_avalon_trace_read                 (abus_slave_0_avalon_trace_read),                   //                                         .read
		.abus_slave_0_avalon_trace_readdata             (abus_slave_0_avalon_trace_readdata),               //                                         .readdata
		.abus_slave_0_avalon_trace_readdatavalid        (abus_slave_0_avalon_trace_readdatavalid),          //                                         .readdatavalid
		.abus_slave_0_avalon_trace_write                (abus_slave_0_avalon_trace_write),                  //                                         .write
		.abus_slave_0_avalon_trace_writedata            (abus_slave_0_avalon_trace_writedata),              //                                         .writedata
		.onchip_trace_mem_s1_address                    (mm_interconnect_1_onchip_trace_mem_s1_address),    //                      onchip_trace_mem_s1.address
		.onchip_trace_mem_s1_write                      (mm_interconnect_1_onchip_trace_mem_s1_write),      //                                         .write
		.onchip_trace_mem_s1_readdata                   (mm_interconnect_1_onchip_trace_mem_s1_readdata),   //                                         .readdata
		.onchip_trace_mem_s1_writedata                  (mm_interconnect_1_onchip_trace_mem_s1_writedata),  //                                         .writedata
		.onchip_trace_mem_s1_byteenable                 (mm_interconnect_1_onchip_trace_mem_s1_byteenable), //                                         .byteenable
		.onchip_trace_mem_s1_chipselect                 (mm_interconnect_1_onchip_trace_mem_s1_chipselect), //                                         .chipselect
		.onchip_trace_mem_s1_clken                      (mm_interconnect_1_onchip_trace_mem_s1_clken)       //                                         .clken
	);

	wasca_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
